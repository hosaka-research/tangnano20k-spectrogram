module nco_rom_4ch_log4943_fs11718 (clock,addr,dataout);
	input clock;
	input [10:0] addr;
	output reg signed [35:0] dataout;
	always @(posedge clock) begin
		case (addr)
			11'h000: dataout<=36'h3c6023c8a;
			11'h001: dataout<=36'h9586d1c2a;
			11'h002: dataout<=36'h7f64bce53;
			11'h003: dataout<=36'h89cf73b6f;
			11'h004: dataout<=36'h3fc864419;
			11'h005: dataout<=36'h9166901ba;
			11'h006: dataout<=36'h7fff3fd00;
			11'h007: dataout<=36'h90a7b0377;
			11'h008: dataout<=36'h4317e4bfa;
			11'h009: dataout<=36'h8db9ce6a6;
			11'h00a: dataout<=36'h7f8a82b2c;
			11'h00b: dataout<=36'h990aacfcf;
			11'h00c: dataout<=36'h464e65427;
			11'h00d: dataout<=36'h8a7f8cb0f;
			11'h00e: dataout<=36'h7e128587a;
			11'h00f: dataout<=36'ha2cc2a112;
			11'h010: dataout<=36'h496ba5c9b;
			11'h011: dataout<=36'h87b7caf15;
			11'h012: dataout<=36'h7ba20848f;
			11'h013: dataout<=36'hadbca77bf;
			11'h014: dataout<=36'h4c6fa6551;
			11'h015: dataout<=36'h8560c92d6;
			11'h016: dataout<=36'h78474af1e;
			11'h017: dataout<=36'hb9ab25439;
			11'h018: dataout<=36'h4f5ae6e46;
			11'h019: dataout<=36'h8378c766a;
			11'h01a: dataout<=36'h740f8d7e6;
			11'h01b: dataout<=36'hc665a36c8;
			11'h01c: dataout<=36'h522ca7773;
			11'h01d: dataout<=36'h81fe459f3;
			11'h01e: dataout<=36'h6f0bcfe9d;
			11'h01f: dataout<=36'hd3ba21f9b;
			11'h020: dataout<=36'h54e5e80d5;
			11'h021: dataout<=36'h80edc3d83;
			11'h022: dataout<=36'h694bd2318;
			11'h023: dataout<=36'he17760ec9;
			11'h024: dataout<=36'h5785e8a67;
			11'h025: dataout<=36'h804582139;
			11'h026: dataout<=36'h62e15451b;
			11'h027: dataout<=36'hef6d20450;
			11'h028: dataout<=36'h5a0d69426;
			11'h029: dataout<=36'h800240526;
			11'h02a: dataout<=36'h5bdc96487;
			11'h02b: dataout<=36'hfd6d2001b;
			11'h02c: dataout<=36'h5c7c69e0d;
			11'h02d: dataout<=36'h8020be962;
			11'h02e: dataout<=36'h545058136;
			11'h02f: dataout<=36'h0b4be0200;
			11'h030: dataout<=36'h5ed32a818;
			11'h031: dataout<=36'h809d3ce01;
			11'h032: dataout<=36'h4c4e19b10;
			11'h033: dataout<=36'h18e0e09c4;
			11'h034: dataout<=36'h6111eb244;
			11'h035: dataout<=36'h81747b314;
			11'h036: dataout<=36'h43e6db202;
			11'h037: dataout<=36'h26062171d;
			11'h038: dataout<=36'h6338ebc8d;
			11'h039: dataout<=36'h82a2b98ad;
			11'h03a: dataout<=36'h3b2c9c5fe;
			11'h03b: dataout<=36'h3299629b4;
			11'h03c: dataout<=36'h65486c6f0;
			11'h03d: dataout<=36'h842437eda;
			11'h03e: dataout<=36'h322f9d6fe;
			11'h03f: dataout<=36'h3e7c24127;
			11'h040: dataout<=36'h6740ad168;
			11'h041: dataout<=36'h85f4765ac;
			11'h042: dataout<=36'h29019e502;
			11'h043: dataout<=36'h4993a5d0b;
			11'h044: dataout<=36'h69222dbf4;
			11'h045: dataout<=36'h881034d2d;
			11'h046: dataout<=36'h1fb15f00c;
			11'h047: dataout<=36'h53c8a7ced;
			11'h048: dataout<=36'h6aed6e691;
			11'h049: dataout<=36'h8a7333566;
			11'h04a: dataout<=36'h164d9f828;
			11'h04b: dataout<=36'h5d07ea056;
			11'h04c: dataout<=36'h6ca22f13a;
			11'h04d: dataout<=36'h8d18f1e69;
			11'h04e: dataout<=36'h0ce71fd60;
			11'h04f: dataout<=36'h6541ec6cd;
			11'h050: dataout<=36'h6e416fbed;
			11'h051: dataout<=36'h8ffd70839;
			11'h052: dataout<=36'h038a1ffca;
			11'h053: dataout<=36'h6c6aeefd6;
			11'h054: dataout<=36'h6fcb706a8;
			11'h055: dataout<=36'h931cef2de;
			11'h056: dataout<=36'hfa435ff7a;
			11'h057: dataout<=36'h727a31af4;
			11'h058: dataout<=36'h714071169;
			11'h059: dataout<=36'h96736de5f;
			11'h05a: dataout<=36'hf11f1fc85;
			11'h05b: dataout<=36'h776af47ae;
			11'h05c: dataout<=36'h72a0b1c2b;
			11'h05d: dataout<=36'h99fc2cac6;
			11'h05e: dataout<=36'he82a1f708;
			11'h05f: dataout<=36'h7b3b3758b;
			11'h060: dataout<=36'h73ed326ef;
			11'h061: dataout<=36'h9db46b80f;
			11'h062: dataout<=36'hdf6bdef21;
			11'h063: dataout<=36'h7debfa419;
			11'h064: dataout<=36'h7525b31b0;
			11'h065: dataout<=36'ha1972a647;
			11'h066: dataout<=36'hd6f09e4ee;
			11'h067: dataout<=36'h7f80bd2e8;
			11'h068: dataout<=36'h764af3c6d;
			11'h069: dataout<=36'ha5a12956b;
			11'h06a: dataout<=36'hcebf9d891;
			11'h06b: dataout<=36'h7fffc018d;
			11'h06c: dataout<=36'h775d74724;
			11'h06d: dataout<=36'ha9ce6857e;
			11'h06e: dataout<=36'hc6e09ca2e;
			11'h06f: dataout<=36'h7f71c2fa6;
			11'h070: dataout<=36'h785d751d4;
			11'h071: dataout<=36'hae1be7682;
			11'h072: dataout<=36'hbf5a1b9e2;
			11'h073: dataout<=36'h7de085cd8;
			11'h074: dataout<=36'h794b75c7a;
			11'h075: dataout<=36'hb285a6877;
			11'h076: dataout<=36'hb832da7d6;
			11'h077: dataout<=36'h7b58c88cb;
			11'h078: dataout<=36'h7a2836714;
			11'h079: dataout<=36'hb707a5b5a;
			11'h07a: dataout<=36'hb16ed9432;
			11'h07b: dataout<=36'h77e74b332;
			11'h07c: dataout<=36'h7af3771a2;
			11'h07d: dataout<=36'hbb9fe4f2f;
			11'h07e: dataout<=36'hab1397f10;
			11'h07f: dataout<=36'h739b4dbc7;
			11'h080: dataout<=36'h7bae37c21;
			11'h081: dataout<=36'hc04a243f0;
			11'h082: dataout<=36'ha523d689d;
			11'h083: dataout<=36'h6e849024b;
			11'h084: dataout<=36'h7c58b8690;
			11'h085: dataout<=36'hc503a399d;
			11'h086: dataout<=36'h9fa2d50fb;
			11'h087: dataout<=36'h68b352688;
			11'h088: dataout<=36'h7cf3790ee;
			11'h089: dataout<=36'hc9c9a3032;
			11'h08a: dataout<=36'h9a925384d;
			11'h08b: dataout<=36'h62389484e;
			11'h08c: dataout<=36'h7d7eb9b3a;
			11'h08d: dataout<=36'hce99627ae;
			11'h08e: dataout<=36'h95f411eb3;
			11'h08f: dataout<=36'h5b2616776;
			11'h090: dataout<=36'h7dfb3a572;
			11'h091: dataout<=36'hd36fe200a;
			11'h092: dataout<=36'h91c890454;
			11'h093: dataout<=36'h538d983df;
			11'h094: dataout<=36'h7e693af95;
			11'h095: dataout<=36'hd84a61944;
			11'h096: dataout<=36'h8e104e951;
			11'h097: dataout<=36'h4b8059d71;
			11'h098: dataout<=36'h7ec8fb9a3;
			11'h099: dataout<=36'hdd2721358;
			11'h09a: dataout<=36'h8acb0cdc5;
			11'h09b: dataout<=36'h43105b419;
			11'h09c: dataout<=36'h7f1afc39b;
			11'h09d: dataout<=36'he203a0e42;
			11'h09e: dataout<=36'h87f88b1d1;
			11'h09f: dataout<=36'h3a4e9c7cb;
			11'h0a0: dataout<=36'h7f5ffcd7a;
			11'h0a1: dataout<=36'he6dca09fa;
			11'h0a2: dataout<=36'h85964959a;
			11'h0a3: dataout<=36'h314c5d880;
			11'h0a4: dataout<=36'h7f97fd742;
			11'h0a5: dataout<=36'hebb1a067d;
			11'h0a6: dataout<=36'h83a387931;
			11'h0a7: dataout<=36'h2819de639;
			11'h0a8: dataout<=36'h7fc37e0f1;
			11'h0a9: dataout<=36'hf07fe03c6;
			11'h0aa: dataout<=36'h821e45cb8;
			11'h0ab: dataout<=36'h1ec6df0fa;
			11'h0ac: dataout<=36'h7fe2fea85;
			11'h0ad: dataout<=36'hf544e01cf;
			11'h0ae: dataout<=36'h8103c404a;
			11'h0af: dataout<=36'h1562df8cd;
			11'h0b0: dataout<=36'h7ff6bf400;
			11'h0b1: dataout<=36'hfa0060092;
			11'h0b2: dataout<=36'h8051823f9;
			11'h0b3: dataout<=36'h0bfc1fdc0;
			11'h0b4: dataout<=36'h7fff7fd60;
			11'h0b5: dataout<=36'hfeb020008;
			11'h0b6: dataout<=36'h8004007df;
			11'h0b7: dataout<=36'h02a05ffe4;
			11'h0b8: dataout<=36'h7ffcc06a2;
			11'h0b9: dataout<=36'h03512002f;
			11'h0ba: dataout<=36'h8019fec19;
			11'h0bb: dataout<=36'hf95cdff4f;
			11'h0bc: dataout<=36'h7ff000fcb;
			11'h0bd: dataout<=36'h07e4e00fb;
			11'h0be: dataout<=36'h808cfd0ac;
			11'h0bf: dataout<=36'hf03d1fc1a;
			11'h0c0: dataout<=36'h7fd9018d8;
			11'h0c1: dataout<=36'h0c686026b;
			11'h0c2: dataout<=36'h815b7b5b3;
			11'h0c3: dataout<=36'he74c9f660;
			11'h0c4: dataout<=36'h7fb8421c8;
			11'h0c5: dataout<=36'h10dae0477;
			11'h0c6: dataout<=36'h828179b3d;
			11'h0c7: dataout<=36'hde951ee3e;
			11'h0c8: dataout<=36'h7f8e02a9b;
			11'h0c9: dataout<=36'h153ae0719;
			11'h0ca: dataout<=36'h83fab815b;
			11'h0cb: dataout<=36'hd6209e3d3;
			11'h0cc: dataout<=36'h7f5a83351;
			11'h0cd: dataout<=36'h1987a0a4c;
			11'h0ce: dataout<=36'h85c43681c;
			11'h0cf: dataout<=36'hcdf71d742;
			11'h0d0: dataout<=36'h7f1e83be9;
			11'h0d1: dataout<=36'h1dc020e07;
			11'h0d2: dataout<=36'h87d834f8b;
			11'h0d3: dataout<=36'hc6205c8ac;
			11'h0d4: dataout<=36'h7eda04464;
			11'h0d5: dataout<=36'h21e3a1247;
			11'h0d6: dataout<=36'h8a33f37b5;
			11'h0d7: dataout<=36'hbea2db835;
			11'h0d8: dataout<=36'h7e8d44cc1;
			11'h0d9: dataout<=36'h25f1a1705;
			11'h0da: dataout<=36'h8cd3720a2;
			11'h0db: dataout<=36'hb784da600;
			11'h0dc: dataout<=36'h7e38c5501;
			11'h0dd: dataout<=36'h29e9a1c3c;
			11'h0de: dataout<=36'h8fb270a5c;
			11'h0df: dataout<=36'hb0cb59233;
			11'h0e0: dataout<=36'h7ddd05d22;
			11'h0e1: dataout<=36'h2dca621e3;
			11'h0e2: dataout<=36'h92cbaf4ec;
			11'h0e3: dataout<=36'haa7a17cf0;
			11'h0e4: dataout<=36'h7d79c6526;
			11'h0e5: dataout<=36'h3193e27f9;
			11'h0e6: dataout<=36'h961d2e058;
			11'h0e7: dataout<=36'ha4951665e;
			11'h0e8: dataout<=36'h7d0fc6d0b;
			11'h0e9: dataout<=36'h354562e75;
			11'h0ea: dataout<=36'h99a1acca7;
			11'h0eb: dataout<=36'h9f1ed4e9f;
			11'h0ec: dataout<=36'h7c9f474d2;
			11'h0ed: dataout<=36'h38dea3551;
			11'h0ee: dataout<=36'h9d54ab9dd;
			11'h0ef: dataout<=36'h9a19935d7;
			11'h0f0: dataout<=36'h7c2847c7c;
			11'h0f1: dataout<=36'h3c5fe3c8b;
			11'h0f2: dataout<=36'ha133ea7fc;
			11'h0f3: dataout<=36'h958651c2a;
			11'h0f4: dataout<=36'h7bab48407;
			11'h0f5: dataout<=36'h3fc7e441a;
			11'h0f6: dataout<=36'ha53a2970a;
			11'h0f7: dataout<=36'h9166501b9;
			11'h0f8: dataout<=36'h7b2888b75;
			11'h0f9: dataout<=36'h4317a4bfb;
			11'h0fa: dataout<=36'ha96468704;
			11'h0fb: dataout<=36'h8db94e6a5;
			11'h0fc: dataout<=36'h7aa0492c4;
			11'h0fd: dataout<=36'h464da5428;
			11'h0fe: dataout<=36'hadaea77f2;
			11'h0ff: dataout<=36'h8a7f8cb0f;
			11'h100: dataout<=36'h7a12c99f7;
			11'h101: dataout<=36'h496b65c9c;
			11'h102: dataout<=36'hb215a69cc;
			11'h103: dataout<=36'h87b78af15;
			11'h104: dataout<=36'h79804a10b;
			11'h105: dataout<=36'h4c6f26552;
			11'h106: dataout<=36'hb695a5c9c;
			11'h107: dataout<=36'h8560892d5;
			11'h108: dataout<=36'h78e90a802;
			11'h109: dataout<=36'h4f5a26e46;
			11'h10a: dataout<=36'hbb2b65058;
			11'h10b: dataout<=36'h83788766b;
			11'h10c: dataout<=36'h784d4aedc;
			11'h10d: dataout<=36'h522c27773;
			11'h10e: dataout<=36'hbfd3e4502;
			11'h10f: dataout<=36'h81fdc59f2;
			11'h110: dataout<=36'h77ad0b599;
			11'h111: dataout<=36'h54e5280d5;
			11'h112: dataout<=36'hc48c63a98;
			11'h113: dataout<=36'h80ed83d84;
			11'h114: dataout<=36'h7708cbc39;
			11'h115: dataout<=36'h578568a68;
			11'h116: dataout<=36'hc95163117;
			11'h117: dataout<=36'h804542138;
			11'h118: dataout<=36'h7660cc2bd;
			11'h119: dataout<=36'h5a0d29426;
			11'h11a: dataout<=36'hce202287a;
			11'h11b: dataout<=36'h8001c0526;
			11'h11c: dataout<=36'h75b50c924;
			11'h11d: dataout<=36'h5c7be9e0c;
			11'h11e: dataout<=36'hd2f5a20c1;
			11'h11f: dataout<=36'h80203e963;
			11'h120: dataout<=36'h7505ccf6f;
			11'h121: dataout<=36'h5ed2aa817;
			11'h122: dataout<=36'hd7d0219e6;
			11'h123: dataout<=36'h809cfce02;
			11'h124: dataout<=36'h74534d59e;
			11'h125: dataout<=36'h61116b243;
			11'h126: dataout<=36'hdcaca13e5;
			11'h127: dataout<=36'h81743b315;
			11'h128: dataout<=36'h739d8dbb2;
			11'h129: dataout<=36'h63386bc8d;
			11'h12a: dataout<=36'he18960eb9;
			11'h12b: dataout<=36'h82a2798ad;
			11'h12c: dataout<=36'h72e50e1aa;
			11'h12d: dataout<=36'h6547ec6ef;
			11'h12e: dataout<=36'he662e0a5e;
			11'h12f: dataout<=36'h8423f7edb;
			11'h130: dataout<=36'h7229ce787;
			11'h131: dataout<=36'h67402d168;
			11'h132: dataout<=36'heb38206ce;
			11'h133: dataout<=36'h85f4765ac;
			11'h134: dataout<=36'h716c0ed4a;
			11'h135: dataout<=36'h69222dbf4;
			11'h136: dataout<=36'hf00720401;
			11'h137: dataout<=36'h881034d2c;
			11'h138: dataout<=36'h70abcf2f1;
			11'h139: dataout<=36'h6aecee690;
			11'h13a: dataout<=36'hf4cd601f9;
			11'h13b: dataout<=36'h8a72f3567;
			11'h13c: dataout<=36'h6fe94f87f;
			11'h13d: dataout<=36'h6ca1ef139;
			11'h13e: dataout<=36'hf989e00aa;
			11'h13f: dataout<=36'h8d18b1e68;
			11'h140: dataout<=36'h6f24cfdf3;
			11'h141: dataout<=36'h6e412fbed;
			11'h142: dataout<=36'hfe3aa000f;
			11'h143: dataout<=36'h8ffd30838;
			11'h144: dataout<=36'h6e5e5034d;
			11'h145: dataout<=36'h6fcaf06a9;
			11'h146: dataout<=36'h02de60025;
			11'h147: dataout<=36'h931caf2dd;
			11'h148: dataout<=36'h6d961088e;
			11'h149: dataout<=36'h713ff1169;
			11'h14a: dataout<=36'h0773600e2;
			11'h14b: dataout<=36'h96732de5f;
			11'h14c: dataout<=36'h6ccc50db6;
			11'h14d: dataout<=36'h72a071c2b;
			11'h14e: dataout<=36'h0bf820241;
			11'h14f: dataout<=36'h99fc2cac4;
			11'h150: dataout<=36'h6c01112c5;
			11'h151: dataout<=36'h73ecb26ee;
			11'h152: dataout<=36'h106c2043e;
			11'h153: dataout<=36'h9db42b810;
			11'h154: dataout<=36'h6b34517bc;
			11'h155: dataout<=36'h7525331af;
			11'h156: dataout<=36'h14cde06d2;
			11'h157: dataout<=36'ha196ea646;
			11'h158: dataout<=36'h6a6651c9b;
			11'h159: dataout<=36'h764a33c6d;
			11'h15a: dataout<=36'h191ca09f8;
			11'h15b: dataout<=36'ha5a0e956a;
			11'h15c: dataout<=36'h699752163;
			11'h15d: dataout<=36'h775cf4724;
			11'h15e: dataout<=36'h1d5760da6;
			11'h15f: dataout<=36'ha9ce6857e;
			11'h160: dataout<=36'h68c752613;
			11'h161: dataout<=36'h785cf51d3;
			11'h162: dataout<=36'h217ce11d9;
			11'h163: dataout<=36'hae1ba7681;
			11'h164: dataout<=36'h67f652aac;
			11'h165: dataout<=36'h794af5c79;
			11'h166: dataout<=36'h258d2168c;
			11'h167: dataout<=36'hb28526875;
			11'h168: dataout<=36'h672492f2f;
			11'h169: dataout<=36'h7a2776714;
			11'h16a: dataout<=36'h298721bb7;
			11'h16b: dataout<=36'hb707a5b5a;
			11'h16c: dataout<=36'h66525339b;
			11'h16d: dataout<=36'h7af2f71a1;
			11'h16e: dataout<=36'h2d6a22153;
			11'h16f: dataout<=36'hbb9fa4f2e;
			11'h170: dataout<=36'h657f537f1;
			11'h171: dataout<=36'h7bad77c20;
			11'h172: dataout<=36'h3135a275f;
			11'h173: dataout<=36'hc049e43ef;
			11'h174: dataout<=36'h64ac13c32;
			11'h175: dataout<=36'h7c587868e;
			11'h176: dataout<=36'h34e9a2dce;
			11'h177: dataout<=36'hc503a399c;
			11'h178: dataout<=36'h63d81405d;
			11'h179: dataout<=36'h7cf2b90ed;
			11'h17a: dataout<=36'h3885634a5;
			11'h17b: dataout<=36'hc9c9a3031;
			11'h17c: dataout<=36'h630414474;
			11'h17d: dataout<=36'h7d7e79b3a;
			11'h17e: dataout<=36'h3c0963bd4;
			11'h17f: dataout<=36'hce99227ac;
			11'h180: dataout<=36'h622fd4876;
			11'h181: dataout<=36'h7dfafa572;
			11'h182: dataout<=36'h3f742435b;
			11'h183: dataout<=36'hd36fa2009;
			11'h184: dataout<=36'h615b94c63;
			11'h185: dataout<=36'h7e68baf94;
			11'h186: dataout<=36'h42c5a4b33;
			11'h187: dataout<=36'hd84a61944;
			11'h188: dataout<=36'h60871503c;
			11'h189: dataout<=36'h7ec83b9a2;
			11'h18a: dataout<=36'h45fe2535a;
			11'h18b: dataout<=36'hdd2721358;
			11'h18c: dataout<=36'h5fb2d5402;
			11'h18d: dataout<=36'h7f1abc399;
			11'h18e: dataout<=36'h491e25bc5;
			11'h18f: dataout<=36'he20360e40;
			11'h190: dataout<=36'h5ede957b5;
			11'h191: dataout<=36'h7f5fbcd79;
			11'h192: dataout<=36'h4c24e6475;
			11'h193: dataout<=36'he6dca09f9;
			11'h194: dataout<=36'h5e0a95b54;
			11'h195: dataout<=36'h7f977d740;
			11'h196: dataout<=36'h4f1226d63;
			11'h197: dataout<=36'hebb1a067d;
			11'h198: dataout<=36'h5d3695ee1;
			11'h199: dataout<=36'h7fc2fe0f0;
			11'h19a: dataout<=36'h51e6e768d;
			11'h19b: dataout<=36'hf07fa03c5;
			11'h19c: dataout<=36'h5c635625b;
			11'h19d: dataout<=36'h7fe27ea83;
			11'h19e: dataout<=36'h54a1e7fe8;
			11'h19f: dataout<=36'hf545201ce;
			11'h1a0: dataout<=36'h5b90165c4;
			11'h1a1: dataout<=36'h7ff67f400;
			11'h1a2: dataout<=36'h574528978;
			11'h1a3: dataout<=36'hfa0060091;
			11'h1a4: dataout<=36'h5abd9691a;
			11'h1a5: dataout<=36'h7ffeffd5e;
			11'h1a6: dataout<=36'h59ce69331;
			11'h1a7: dataout<=36'hfeafe0007;
			11'h1a8: dataout<=36'h59eb56c5f;
			11'h1a9: dataout<=36'h7ffc006a3;
			11'h1aa: dataout<=36'h5c3fa9d16;
			11'h1ab: dataout<=36'h0351e002d;
			11'h1ac: dataout<=36'h5919d6f94;
			11'h1ad: dataout<=36'h7fefc0fcd;
			11'h1ae: dataout<=36'h5e99aa71d;
			11'h1af: dataout<=36'h07e5600fa;
			11'h1b0: dataout<=36'h5848d72b7;
			11'h1b1: dataout<=36'h7fd8818da;
			11'h1b2: dataout<=36'h60da6b147;
			11'h1b3: dataout<=36'h0c68e026a;
			11'h1b4: dataout<=36'h5778975c9;
			11'h1b5: dataout<=36'h7fb7821c8;
			11'h1b6: dataout<=36'h63032bb8c;
			11'h1b7: dataout<=36'h10db20476;
			11'h1b8: dataout<=36'h56a9178cc;
			11'h1b9: dataout<=36'h7f8d82a9c;
			11'h1ba: dataout<=36'h65156c5ec;
			11'h1bb: dataout<=36'h153b20718;
			11'h1bc: dataout<=36'h55da57bbf;
			11'h1bd: dataout<=36'h7f5a83352;
			11'h1be: dataout<=36'h67106d062;
			11'h1bf: dataout<=36'h1987e0a4a;
			11'h1c0: dataout<=36'h550c57ea1;
			11'h1c1: dataout<=36'h7f1e03be9;
			11'h1c2: dataout<=36'h68f32daec;
			11'h1c3: dataout<=36'h1dc0a0e06;
			11'h1c4: dataout<=36'h543f18175;
			11'h1c5: dataout<=36'h7ed984465;
			11'h1c6: dataout<=36'h6ac0ee588;
			11'h1c7: dataout<=36'h21e461247;
			11'h1c8: dataout<=36'h5372d8439;
			11'h1c9: dataout<=36'h7e8cc4cc1;
			11'h1ca: dataout<=36'h6c77af02f;
			11'h1cb: dataout<=36'h25f261705;
			11'h1cc: dataout<=36'h52a7586ef;
			11'h1cd: dataout<=36'h7e3845502;
			11'h1ce: dataout<=36'h6e192fae3;
			11'h1cf: dataout<=36'h29ea21c3b;
			11'h1d0: dataout<=36'h51dd18996;
			11'h1d1: dataout<=36'h7ddc85d22;
			11'h1d2: dataout<=36'h6fa4f059b;
			11'h1d3: dataout<=36'h2dcae21e3;
			11'h1d4: dataout<=36'h511398c2f;
			11'h1d5: dataout<=36'h7d7946526;
			11'h1d6: dataout<=36'h711bf105c;
			11'h1d7: dataout<=36'h3194627f8;
			11'h1d8: dataout<=36'h504b18eba;
			11'h1d9: dataout<=36'h7d0f46d0b;
			11'h1da: dataout<=36'h727e71b1f;
			11'h1db: dataout<=36'h3545e2e74;
			11'h1dc: dataout<=36'h4f83d9138;
			11'h1dd: dataout<=36'h7c9f074d3;
			11'h1de: dataout<=36'h73cd325e1;
			11'h1df: dataout<=36'h38df63551;
			11'h1e0: dataout<=36'h4ebd593a7;
			11'h1e1: dataout<=36'h7c2787c7c;
			11'h1e2: dataout<=36'h7506f30a4;
			11'h1e3: dataout<=36'h3c6063c8a;
			11'h1e4: dataout<=36'h4df85960a;
			11'h1e5: dataout<=36'h7bab08407;
			11'h1e6: dataout<=36'h762e73b60;
			11'h1e7: dataout<=36'h3fc8a4419;
			11'h1e8: dataout<=36'h4d3419860;
			11'h1e9: dataout<=36'h7b2808b76;
			11'h1ea: dataout<=36'h7742b461b;
			11'h1eb: dataout<=36'h431824bfa;
			11'h1ec: dataout<=36'h4c7159aa9;
			11'h1ed: dataout<=36'h7aa0092c5;
			11'h1ee: dataout<=36'h7844b50c9;
			11'h1ef: dataout<=36'h464ea5427;
			11'h1f0: dataout<=36'h4baf99ce5;
			11'h1f1: dataout<=36'h7a12499f6;
			11'h1f2: dataout<=36'h7933f5b6f;
			11'h1f3: dataout<=36'h496be5c9b;
			11'h1f4: dataout<=36'h4aef19f16;
			11'h1f5: dataout<=36'h79800a10c;
			11'h1f6: dataout<=36'h7a12b660c;
			11'h1f7: dataout<=36'h4c6fe6551;
			11'h1f8: dataout<=36'h4a2f9a13a;
			11'h1f9: dataout<=36'h78e88a803;
			11'h1fa: dataout<=36'h7adf7709b;
			11'h1fb: dataout<=36'h4f5b26e46;
			11'h1fc: dataout<=36'h49719a353;
			11'h1fd: dataout<=36'h784ccaedd;
			11'h1fe: dataout<=36'h7b9bf7b1b;
			11'h1ff: dataout<=36'h522ce7773;
			11'h200: dataout<=36'h48b4da560;
			11'h201: dataout<=36'h77accb599;
			11'h202: dataout<=36'h7c47f858b;
			11'h203: dataout<=36'h54e6280d5;
			11'h204: dataout<=36'h47f91a762;
			11'h205: dataout<=36'h77084bc3a;
			11'h206: dataout<=36'h7ce438fec;
			11'h207: dataout<=36'h578628a67;
			11'h208: dataout<=36'h473eda959;
			11'h209: dataout<=36'h76604c2bd;
			11'h20a: dataout<=36'h7d70f9a39;
			11'h20b: dataout<=36'h5a0da9426;
			11'h20c: dataout<=36'h4685dab45;
			11'h20d: dataout<=36'h75b44c924;
			11'h20e: dataout<=36'h7dee7a473;
			11'h20f: dataout<=36'h5c7ca9e0d;
			11'h210: dataout<=36'h45ce1ad27;
			11'h211: dataout<=36'h75050cf70;
			11'h212: dataout<=36'h7e5dfae9a;
			11'h213: dataout<=36'h5ed36a818;
			11'h214: dataout<=36'h4517daefe;
			11'h215: dataout<=36'h7452cd59e;
			11'h216: dataout<=36'h7ebf3b8a8;
			11'h217: dataout<=36'h61122b244;
			11'h218: dataout<=36'h4462db0cb;
			11'h219: dataout<=36'h739d0dbb2;
			11'h21a: dataout<=36'h7f12bc2a2;
			11'h21b: dataout<=36'h63392bc8d;
			11'h21c: dataout<=36'h43af1b28e;
			11'h21d: dataout<=36'h72e48e1aa;
			11'h21e: dataout<=36'h7f58fcc84;
			11'h21f: dataout<=36'h6548ac6f0;
			11'h220: dataout<=36'h42fcdb447;
			11'h221: dataout<=36'h72294e786;
			11'h222: dataout<=36'h7f91fd64d;
			11'h223: dataout<=36'h6740ed168;
			11'h224: dataout<=36'h424bdb5f7;
			11'h225: dataout<=36'h716b8ed49;
			11'h226: dataout<=36'h7fbefdffe;
			11'h227: dataout<=36'h69226dbf4;
			11'h228: dataout<=36'h419c1b79e;
			11'h229: dataout<=36'h70ab4f2f3;
			11'h22a: dataout<=36'h7fdffe998;
			11'h22b: dataout<=36'h6aedae691;
			11'h22c: dataout<=36'h40eddb93b;
			11'h22d: dataout<=36'h6fe8cf880;
			11'h22e: dataout<=36'h7ff4bf315;
			11'h22f: dataout<=36'h6ca26f13a;
			11'h230: dataout<=36'h40411bacf;
			11'h231: dataout<=36'h6f248fdf3;
			11'h232: dataout<=36'h7ffe7fc76;
			11'h233: dataout<=36'h6e41afbed;
			11'h234: dataout<=36'h3f959bc5a;
			11'h235: dataout<=36'h6e5dd034d;
			11'h236: dataout<=36'h7ffc805bd;
			11'h237: dataout<=36'h6fcbb06a8;
			11'h238: dataout<=36'h3eeb5bddd;
			11'h239: dataout<=36'h6d959088f;
			11'h23a: dataout<=36'h7ff0c0eea;
			11'h23b: dataout<=36'h7140b1169;
			11'h23c: dataout<=36'h3e42dbf57;
			11'h23d: dataout<=36'h6ccc10db5;
			11'h23e: dataout<=36'h7fdb017f6;
			11'h23f: dataout<=36'h72a0f1c2b;
			11'h240: dataout<=36'h3d9b5c0c9;
			11'h241: dataout<=36'h6c00512c5;
			11'h242: dataout<=36'h7fba820eb;
			11'h243: dataout<=36'h73ed726ef;
			11'h244: dataout<=36'h3cf59c233;
			11'h245: dataout<=36'h6b34117bc;
			11'h246: dataout<=36'h7f91c29bf;
			11'h247: dataout<=36'h7525f31b0;
			11'h248: dataout<=36'h3c511c395;
			11'h249: dataout<=36'h6a6611c9b;
			11'h24a: dataout<=36'h7f5f43278;
			11'h24b: dataout<=36'h764b33c6d;
			11'h24c: dataout<=36'h3baddc4f0;
			11'h24d: dataout<=36'h699712164;
			11'h24e: dataout<=36'h7f2443b15;
			11'h24f: dataout<=36'h775db4724;
			11'h250: dataout<=36'h3b0c1c642;
			11'h251: dataout<=36'h68c6d2613;
			11'h252: dataout<=36'h7ee004392;
			11'h253: dataout<=36'h785db51d4;
			11'h254: dataout<=36'h3a6bdc78e;
			11'h255: dataout<=36'h67f652aad;
			11'h256: dataout<=36'h7e94c4bf2;
			11'h257: dataout<=36'h794bb5c7a;
			11'h258: dataout<=36'h39ccdc8d2;
			11'h259: dataout<=36'h672452f30;
			11'h25a: dataout<=36'h7e4105436;
			11'h25b: dataout<=36'h7a2876714;
			11'h25c: dataout<=36'h392f5ca0e;
			11'h25d: dataout<=36'h6651d339a;
			11'h25e: dataout<=36'h7de545c58;
			11'h25f: dataout<=36'h7af3b71a2;
			11'h260: dataout<=36'h38931cb44;
			11'h261: dataout<=36'h657ed37f1;
			11'h262: dataout<=36'h7d82c645f;
			11'h263: dataout<=36'h7bae77c21;
			11'h264: dataout<=36'h37f85cc73;
			11'h265: dataout<=36'h64ab93c32;
			11'h266: dataout<=36'h7d1986c48;
			11'h267: dataout<=36'h7c58f8690;
			11'h268: dataout<=36'h375edcd9c;
			11'h269: dataout<=36'h63d79405f;
			11'h26a: dataout<=36'h7ca9c7414;
			11'h26b: dataout<=36'h7cf3b90ee;
			11'h26c: dataout<=36'h36c71cebd;
			11'h26d: dataout<=36'h6303d4473;
			11'h26e: dataout<=36'h7c3387bbd;
			11'h26f: dataout<=36'h7d7ef9b3a;
			11'h270: dataout<=36'h36305cfd9;
			11'h271: dataout<=36'h622f94876;
			11'h272: dataout<=36'h7bb74834d;
			11'h273: dataout<=36'h7dfb7a572;
			11'h274: dataout<=36'h359b1d0ee;
			11'h275: dataout<=36'h615b14c63;
			11'h276: dataout<=36'h7b34c8abd;
			11'h277: dataout<=36'h7e697af95;
			11'h278: dataout<=36'h35075d1fd;
			11'h279: dataout<=36'h6086d503d;
			11'h27a: dataout<=36'h7aad89210;
			11'h27b: dataout<=36'h7ec93b9a3;
			11'h27c: dataout<=36'h3474dd306;
			11'h27d: dataout<=36'h5fb295402;
			11'h27e: dataout<=36'h7a2089944;
			11'h27f: dataout<=36'h7f1b3c39b;
			11'h280: dataout<=36'h33e39d409;
			11'h281: dataout<=36'h5ede157b5;
			11'h282: dataout<=36'h798e0a05d;
			11'h283: dataout<=36'h7f603cd7a;
			11'h284: dataout<=36'h3353dd506;
			11'h285: dataout<=36'h5e09d5b54;
			11'h286: dataout<=36'h78f70a756;
			11'h287: dataout<=36'h7f983d742;
			11'h288: dataout<=36'h32c59d5fe;
			11'h289: dataout<=36'h5d3695ee0;
			11'h28a: dataout<=36'h785c0ae31;
			11'h28b: dataout<=36'h7fc3be0f1;
			11'h28c: dataout<=36'h32385d6f0;
			11'h28d: dataout<=36'h5c629625b;
			11'h28e: dataout<=36'h77bbcb4f3;
			11'h28f: dataout<=36'h7fe33ea85;
			11'h290: dataout<=36'h31ac9d7dd;
			11'h291: dataout<=36'h5b8f965c4;
			11'h292: dataout<=36'h77180bb96;
			11'h293: dataout<=36'h7ff6ff400;
			11'h294: dataout<=36'h31225d8c5;
			11'h295: dataout<=36'h5abd5691b;
			11'h296: dataout<=36'h7670cc21c;
			11'h297: dataout<=36'h7fffbfd60;
			11'h298: dataout<=36'h30995d9a7;
			11'h299: dataout<=36'h59eb16c5f;
			11'h29a: dataout<=36'h75c54c885;
			11'h29b: dataout<=36'h7ffd006a3;
			11'h29c: dataout<=36'h30119da85;
			11'h29d: dataout<=36'h591996f94;
			11'h29e: dataout<=36'h75168ced4;
			11'h29f: dataout<=36'h7ff040fcc;
			11'h2a0: dataout<=36'h2f8b1db5d;
			11'h2a1: dataout<=36'h5848972b7;
			11'h2a2: dataout<=36'h74640d506;
			11'h2a3: dataout<=36'h7fd9418d9;
			11'h2a4: dataout<=36'h2f061dc31;
			11'h2a5: dataout<=36'h5778575ca;
			11'h2a6: dataout<=36'h73aecdb1c;
			11'h2a7: dataout<=36'h7fb8821c9;
			11'h2a8: dataout<=36'h2e825dd00;
			11'h2a9: dataout<=36'h56a9178cc;
			11'h2aa: dataout<=36'h72f6ce116;
			11'h2ab: dataout<=36'h7f8e42a9c;
			11'h2ac: dataout<=36'h2dff9ddca;
			11'h2ad: dataout<=36'h55d997bbf;
			11'h2ae: dataout<=36'h723b0e6f8;
			11'h2af: dataout<=36'h7f5ac3352;
			11'h2b0: dataout<=36'h2d7e9de90;
			11'h2b1: dataout<=36'h550c17ea1;
			11'h2b2: dataout<=36'h717e0ecba;
			11'h2b3: dataout<=36'h7f1ec3bea;
			11'h2b4: dataout<=36'h2cfe9df51;
			11'h2b5: dataout<=36'h543ed8174;
			11'h2b6: dataout<=36'h70bdcf264;
			11'h2b7: dataout<=36'h7eda44465;
			11'h2b8: dataout<=36'h2c7fde00e;
			11'h2b9: dataout<=36'h537258439;
			11'h2ba: dataout<=36'h6ffb8f7f5;
			11'h2bb: dataout<=36'h7e8d84cc2;
			11'h2bc: dataout<=36'h2c029e0c7;
			11'h2bd: dataout<=36'h52a7186ef;
			11'h2be: dataout<=36'h6f374fd6c;
			11'h2bf: dataout<=36'h7e3905502;
			11'h2c0: dataout<=36'h2b865e17c;
			11'h2c1: dataout<=36'h51dc98997;
			11'h2c2: dataout<=36'h6e71102ca;
			11'h2c3: dataout<=36'h7ddd45d23;
			11'h2c4: dataout<=36'h2b0b5e22c;
			11'h2c5: dataout<=36'h5112d8c2f;
			11'h2c6: dataout<=36'h6da89080c;
			11'h2c7: dataout<=36'h7d7a06527;
			11'h2c8: dataout<=36'h2a91de2d9;
			11'h2c9: dataout<=36'h504ad8eba;
			11'h2ca: dataout<=36'h6cdf90d36;
			11'h2cb: dataout<=36'h7d1006d0c;
			11'h2cc: dataout<=36'h2a195e382;
			11'h2cd: dataout<=36'h4f8359138;
			11'h2ce: dataout<=36'h6c1411249;
			11'h2cf: dataout<=36'h7c9f874d3;
			11'h2d0: dataout<=36'h29a21e427;
			11'h2d1: dataout<=36'h4ebcd93a8;
			11'h2d2: dataout<=36'h6b4751743;
			11'h2d3: dataout<=36'h7c2887c7d;
			11'h2d4: dataout<=36'h292c1e4c8;
			11'h2d5: dataout<=36'h4df79960a;
			11'h2d6: dataout<=36'h6a7951c23;
			11'h2d7: dataout<=36'h7bab88408;
			11'h2d8: dataout<=36'h28b75e566;
			11'h2d9: dataout<=36'h4d3399860;
			11'h2da: dataout<=36'h69aa920ee;
			11'h2db: dataout<=36'h7b28c8b76;
			11'h2dc: dataout<=36'h2843de600;
			11'h2dd: dataout<=36'h4c70d9aa8;
			11'h2de: dataout<=36'h68dad259e;
			11'h2df: dataout<=36'h7aa0892c5;
			11'h2e0: dataout<=36'h27d15e697;
			11'h2e1: dataout<=36'h4baf19ce6;
			11'h2e2: dataout<=36'h680a12a3c;
			11'h2e3: dataout<=36'h7a13099f8;
			11'h2e4: dataout<=36'h27601e72a;
			11'h2e5: dataout<=36'h4aee59f15;
			11'h2e6: dataout<=36'h673812ebf;
			11'h2e7: dataout<=36'h79808a10c;
			11'h2e8: dataout<=36'h26f01e7ba;
			11'h2e9: dataout<=36'h4a2f1a13a;
			11'h2ea: dataout<=36'h6665d332e;
			11'h2eb: dataout<=36'h78e94a803;
			11'h2ec: dataout<=36'h26815e847;
			11'h2ed: dataout<=36'h49715a353;
			11'h2ee: dataout<=36'h659353786;
			11'h2ef: dataout<=36'h784d8aedd;
			11'h2f0: dataout<=36'h26139e8d1;
			11'h2f1: dataout<=36'h48b49a561;
			11'h2f2: dataout<=36'h64c053bca;
			11'h2f3: dataout<=36'h77ad4b59a;
			11'h2f4: dataout<=36'h25a6de957;
			11'h2f5: dataout<=36'h47f89a762;
			11'h2f6: dataout<=36'h63ebd3ff6;
			11'h2f7: dataout<=36'h77090bc3a;
			11'h2f8: dataout<=36'h253b9e9db;
			11'h2f9: dataout<=36'h473eda959;
			11'h2fa: dataout<=36'h63189440e;
			11'h2fb: dataout<=36'h76610c2be;
			11'h2fc: dataout<=36'h24d11ea5b;
			11'h2fd: dataout<=36'h46855ab45;
			11'h2fe: dataout<=36'h624394812;
			11'h2ff: dataout<=36'h75b54c925;
			11'h300: dataout<=36'h2467dead9;
			11'h301: dataout<=36'h45cddad27;
			11'h302: dataout<=36'h616f94c02;
			11'h303: dataout<=36'h75060cf70;
			11'h304: dataout<=36'h23ffdeb54;
			11'h305: dataout<=36'h45179aefe;
			11'h306: dataout<=36'h609b54fdd;
			11'h307: dataout<=36'h74538d59f;
			11'h308: dataout<=36'h2398debcc;
			11'h309: dataout<=36'h44629b0cb;
			11'h30a: dataout<=36'h5fc7153a5;
			11'h30b: dataout<=36'h739dcdbb3;
			11'h30c: dataout<=36'h2332dec41;
			11'h30d: dataout<=36'h43aedb28e;
			11'h30e: dataout<=36'h5ef295759;
			11'h30f: dataout<=36'h72e54e1ab;
			11'h310: dataout<=36'h22ce1ecb4;
			11'h311: dataout<=36'h42fc9b447;
			11'h312: dataout<=36'h5e1ed5afa;
			11'h313: dataout<=36'h722a0e788;
			11'h314: dataout<=36'h226a1ed24;
			11'h315: dataout<=36'h424b5b5f7;
			11'h316: dataout<=36'h5d4a95e89;
			11'h317: dataout<=36'h716c4ed4b;
			11'h318: dataout<=36'h22079ed91;
			11'h319: dataout<=36'h419c1b79c;
			11'h31a: dataout<=36'h5c7756203;
			11'h31b: dataout<=36'h70ac0f2f2;
			11'h31c: dataout<=36'h21a5dedfc;
			11'h31d: dataout<=36'h40ed9b939;
			11'h31e: dataout<=36'h5ba3d656d;
			11'h31f: dataout<=36'h6fe98f880;
			11'h320: dataout<=36'h21451ee65;
			11'h321: dataout<=36'h40409bace;
			11'h322: dataout<=36'h5ad1168c7;
			11'h323: dataout<=36'h6f250fdf4;
			11'h324: dataout<=36'h20e59eecb;
			11'h325: dataout<=36'h3f955bc59;
			11'h326: dataout<=36'h59ff56c0d;
			11'h327: dataout<=36'h6e5e9034e;
			11'h328: dataout<=36'h20871ef30;
			11'h329: dataout<=36'h3eeb5bddd;
			11'h32a: dataout<=36'h592e16f44;
			11'h32b: dataout<=36'h6d965088f;
			11'h32c: dataout<=36'h20295ef91;
			11'h32d: dataout<=36'h3e425bf57;
			11'h32e: dataout<=36'h585c97269;
			11'h32f: dataout<=36'h6ccc90db7;
			11'h330: dataout<=36'h1fccdeff1;
			11'h331: dataout<=36'h3d9b1c0c9;
			11'h332: dataout<=36'h578c5757d;
			11'h333: dataout<=36'h6c01512c6;
			11'h334: dataout<=36'h1f715f04e;
			11'h335: dataout<=36'h3cf55c232;
			11'h336: dataout<=36'h56bcd7880;
			11'h337: dataout<=36'h6b34917bd;
			11'h338: dataout<=36'h1f169f0a9;
			11'h339: dataout<=36'h3c505c394;
			11'h33a: dataout<=36'h55ed57b74;
			11'h33b: dataout<=36'h6a6691c9c;
			11'h33c: dataout<=36'h1ebd1f103;
			11'h33d: dataout<=36'h3bad9c4f0;
			11'h33e: dataout<=36'h551fd7e5a;
			11'h33f: dataout<=36'h699792164;
			11'h340: dataout<=36'h1e645f15a;
			11'h341: dataout<=36'h3b0b9c642;
			11'h342: dataout<=36'h54521812f;
			11'h343: dataout<=36'h68c792614;
			11'h344: dataout<=36'h1e0cdf1af;
			11'h345: dataout<=36'h3a6b9c78d;
			11'h346: dataout<=36'h5386583f4;
			11'h347: dataout<=36'h67f692aad;
			11'h348: dataout<=36'h1db61f202;
			11'h349: dataout<=36'h39cc9c8d0;
			11'h34a: dataout<=36'h52ba986aa;
			11'h34b: dataout<=36'h6724d2f30;
			11'h34c: dataout<=36'h1d605f254;
			11'h34d: dataout<=36'h392f1ca0e;
			11'h34e: dataout<=36'h51f058954;
			11'h34f: dataout<=36'h66529339c;
			11'h350: dataout<=36'h1d0b5f2a3;
			11'h351: dataout<=36'h38929cb43;
			11'h352: dataout<=36'h512618bee;
			11'h353: dataout<=36'h657f937f2;
			11'h354: dataout<=36'h1cb75f2f1;
			11'h355: dataout<=36'h37f7dcc73;
			11'h356: dataout<=36'h505d98e7b;
			11'h357: dataout<=36'h64ac53c33;
			11'h358: dataout<=36'h1c645f33d;
			11'h359: dataout<=36'h375e5cd9b;
			11'h35a: dataout<=36'h4f96190fa;
			11'h35b: dataout<=36'h63d85405e;
			11'h35c: dataout<=36'h1c125f387;
			11'h35d: dataout<=36'h36c69cebc;
			11'h35e: dataout<=36'h4ed019369;
			11'h35f: dataout<=36'h630454475;
			11'h360: dataout<=36'h1bc11f3d0;
			11'h361: dataout<=36'h36301cfd8;
			11'h362: dataout<=36'h4e0ad95ce;
			11'h363: dataout<=36'h623014877;
			11'h364: dataout<=36'h1b70df417;
			11'h365: dataout<=36'h359add0ed;
			11'h366: dataout<=36'h4d4699825;
			11'h367: dataout<=36'h615bd4c64;
			11'h368: dataout<=36'h1b215f45c;
			11'h369: dataout<=36'h3506dd1fc;
			11'h36a: dataout<=36'h4c8399a6f;
			11'h36b: dataout<=36'h60875503d;
			11'h36c: dataout<=36'h1ad2df4a0;
			11'h36d: dataout<=36'h34749d305;
			11'h36e: dataout<=36'h4bc1d9cad;
			11'h36f: dataout<=36'h5fb315403;
			11'h370: dataout<=36'h1a851f4e2;
			11'h371: dataout<=36'h33e35d408;
			11'h372: dataout<=36'h4b0119ede;
			11'h373: dataout<=36'h5eded57b6;
			11'h374: dataout<=36'h1a381f523;
			11'h375: dataout<=36'h33535d506;
			11'h376: dataout<=36'h4a415a105;
			11'h377: dataout<=36'h5e0ad5b55;
			11'h378: dataout<=36'h19ec1f562;
			11'h379: dataout<=36'h32c51d5fd;
			11'h37a: dataout<=36'h49835a31e;
			11'h37b: dataout<=36'h5d36d5ee2;
			11'h37c: dataout<=36'h19a0df5a0;
			11'h37d: dataout<=36'h3237dd6f0;
			11'h37e: dataout<=36'h48c61a52d;
			11'h37f: dataout<=36'h5c639625c;
			11'h380: dataout<=36'h19569f5dd;
			11'h381: dataout<=36'h31ac5d7de;
			11'h382: dataout<=36'h480ada732;
			11'h383: dataout<=36'h5b90565c5;
			11'h384: dataout<=36'h190d1f618;
			11'h385: dataout<=36'h31221d8c5;
			11'h386: dataout<=36'h47509a929;
			11'h387: dataout<=36'h5abdd691b;
			11'h388: dataout<=36'h18c45f651;
			11'h389: dataout<=36'h3098dd9a6;
			11'h38a: dataout<=36'h46971ab14;
			11'h38b: dataout<=36'h59eb96c60;
			11'h38c: dataout<=36'h187c5f68a;
			11'h38d: dataout<=36'h30111da85;
			11'h38e: dataout<=36'h45df5acf9;
			11'h38f: dataout<=36'h591a16f95;
			11'h390: dataout<=36'h18355f6c1;
			11'h391: dataout<=36'h2f8addb5d;
			11'h392: dataout<=36'h45291aed0;
			11'h393: dataout<=36'h5849172b8;
			11'h394: dataout<=36'h17eedf6f7;
			11'h395: dataout<=36'h2f059dc31;
			11'h396: dataout<=36'h44739b09f;
			11'h397: dataout<=36'h5778d75ca;
			11'h398: dataout<=36'h17a95f72b;
			11'h399: dataout<=36'h2e81ddcff;
			11'h39a: dataout<=36'h43bfdb261;
			11'h39b: dataout<=36'h56a9578cd;
			11'h39c: dataout<=36'h17649f75f;
			11'h39d: dataout<=36'h2dff5ddca;
			11'h39e: dataout<=36'h430d5b41d;
			11'h39f: dataout<=36'h55da97bc0;
			11'h3a0: dataout<=36'h17209f791;
			11'h3a1: dataout<=36'h2d7e1de8f;
			11'h3a2: dataout<=36'h425c5b5cc;
			11'h3a3: dataout<=36'h550c97ea2;
			11'h3a4: dataout<=36'h16dd5f7c2;
			11'h3a5: dataout<=36'h2cfe5df50;
			11'h3a6: dataout<=36'h41ac9b773;
			11'h3a7: dataout<=36'h543f58176;
			11'h3a8: dataout<=36'h169adf7f2;
			11'h3a9: dataout<=36'h2c7f9e00d;
			11'h3aa: dataout<=36'h40fe5b911;
			11'h3ab: dataout<=36'h53731843a;
			11'h3ac: dataout<=36'h16591f821;
			11'h3ad: dataout<=36'h2c025e0c6;
			11'h3ae: dataout<=36'h40515baa6;
			11'h3af: dataout<=36'h52a7986f0;
			11'h3b0: dataout<=36'h1617df84f;
			11'h3b1: dataout<=36'h2b85de17b;
			11'h3b2: dataout<=36'h3fa55bc33;
			11'h3b3: dataout<=36'h51dd58997;
			11'h3b4: dataout<=36'h15d79f87c;
			11'h3b5: dataout<=36'h2b0b1e22c;
			11'h3b6: dataout<=36'h3efb5bdb7;
			11'h3b7: dataout<=36'h5113d8c30;
			11'h3b8: dataout<=36'h15981f8a8;
			11'h3b9: dataout<=36'h2a919e2d9;
			11'h3ba: dataout<=36'h3e52dbf32;
			11'h3bb: dataout<=36'h504b58ebb;
			11'h3bc: dataout<=36'h15591f8d2;
			11'h3bd: dataout<=36'h2a191e380;
			11'h3be: dataout<=36'h3daadc0a3;
			11'h3bf: dataout<=36'h4f8419139;
			11'h3c0: dataout<=36'h151adf8fc;
			11'h3c1: dataout<=36'h29a19e426;
			11'h3c2: dataout<=36'h3d049c20f;
			11'h3c3: dataout<=36'h4ebd993a8;
			11'h3c4: dataout<=36'h14dd5f925;
			11'h3c5: dataout<=36'h292bde4c7;
			11'h3c6: dataout<=36'h3c601c371;
			11'h3c7: dataout<=36'h4df89960b;
			11'h3c8: dataout<=36'h14a09f94d;
			11'h3c9: dataout<=36'h28b71e565;
			11'h3ca: dataout<=36'h3bbd1c4cd;
			11'h3cb: dataout<=36'h4d3459861;
			11'h3cc: dataout<=36'h14645f974;
			11'h3cd: dataout<=36'h28435e5ff;
			11'h3ce: dataout<=36'h3b1adc620;
			11'h3cf: dataout<=36'h4c7199aaa;
			11'h3d0: dataout<=36'h14291f99a;
			11'h3d1: dataout<=36'h27d15e695;
			11'h3d2: dataout<=36'h3a7adc76b;
			11'h3d3: dataout<=36'h4bafd9ce6;
			11'h3d4: dataout<=36'h13ee1f9c0;
			11'h3d5: dataout<=36'h275f9e72a;
			11'h3d6: dataout<=36'h39db5c8b2;
			11'h3d7: dataout<=36'h4aef59f17;
			11'h3d8: dataout<=36'h13b41f9e4;
			11'h3d9: dataout<=36'h26efde7b9;
			11'h3da: dataout<=36'h393ddc9ee;
			11'h3db: dataout<=36'h4a2fda13b;
			11'h3dc: dataout<=36'h137a9fa08;
			11'h3dd: dataout<=36'h26811e847;
			11'h3de: dataout<=36'h38a1dcb26;
			11'h3df: dataout<=36'h4971da354;
			11'h3e0: dataout<=36'h1341dfa2b;
			11'h3e1: dataout<=36'h26135e8d1;
			11'h3e2: dataout<=36'h38071cc56;
			11'h3e3: dataout<=36'h48b51a561;
			11'h3e4: dataout<=36'h13099fa4d;
			11'h3e5: dataout<=36'h25a6de957;
			11'h3e6: dataout<=36'h376d9cd7f;
			11'h3e7: dataout<=36'h47f95a763;
			11'h3e8: dataout<=36'h12d21fa6e;
			11'h3e9: dataout<=36'h253b5e9da;
			11'h3ea: dataout<=36'h36d55cea0;
			11'h3eb: dataout<=36'h473f1a95a;
			11'h3ec: dataout<=36'h129b1fa8e;
			11'h3ed: dataout<=36'h24d0dea5a;
			11'h3ee: dataout<=36'h363e5cfbb;
			11'h3ef: dataout<=36'h46861ab46;
			11'h3f0: dataout<=36'h12649faae;
			11'h3f1: dataout<=36'h24675ead8;
			11'h3f2: dataout<=36'h35a89d0d2;
			11'h3f3: dataout<=36'h45ce5ad28;
			11'h3f4: dataout<=36'h122f1facd;
			11'h3f5: dataout<=36'h23ff9eb53;
			11'h3f6: dataout<=36'h35151d1e1;
			11'h3f7: dataout<=36'h45181aeff;
			11'h3f8: dataout<=36'h11f9dfaeb;
			11'h3f9: dataout<=36'h23985ebca;
			11'h3fa: dataout<=36'h34821d2ea;
			11'h3fb: dataout<=36'h44631b0cc;
			11'h3fc: dataout<=36'h11c55fb09;
			11'h3fd: dataout<=36'h23329ec40;
			11'h3fe: dataout<=36'h33f11d3ee;
			11'h3ff: dataout<=36'h43af5b28f;
			11'h400: dataout<=36'h11915fb26;
			11'h401: dataout<=36'h22cd9ecb3;
			11'h402: dataout<=36'h33611d4ed;
			11'h403: dataout<=36'h42fd1b448;
			11'h404: dataout<=36'h115e1fb42;
			11'h405: dataout<=36'h2269ded23;
			11'h406: dataout<=36'h32d29d5e5;
			11'h407: dataout<=36'h424c1b5f8;
			11'h408: dataout<=36'h112b5fb5e;
			11'h409: dataout<=36'h22071ed91;
			11'h40a: dataout<=36'h32455d6d8;
			11'h40b: dataout<=36'h419c5b79f;
			11'h40c: dataout<=36'h10f91fb79;
			11'h40d: dataout<=36'h21a55edfc;
			11'h40e: dataout<=36'h31b99d7c6;
			11'h40f: dataout<=36'h40ee1b93c;
			11'h410: dataout<=36'h10c79fb93;
			11'h411: dataout<=36'h21451ee64;
			11'h412: dataout<=36'h312f5d8ac;
			11'h413: dataout<=36'h40415bad0;
			11'h414: dataout<=36'h10965fbad;
			11'h415: dataout<=36'h20e51eecb;
			11'h416: dataout<=36'h30a59d990;
			11'h417: dataout<=36'h3f95dbc5b;
			11'h418: dataout<=36'h1065dfbc6;
			11'h419: dataout<=36'h20865ef2e;
			11'h41a: dataout<=36'h301d9da6d;
			11'h41b: dataout<=36'h3eeb9bdde;
			11'h41c: dataout<=36'h10361fbdf;
			11'h41d: dataout<=36'h20295ef91;
			11'h41e: dataout<=36'h2f97ddb47;
			11'h41f: dataout<=36'h3e431bf58;
			11'h420: dataout<=36'h10069fbf7;
			11'h421: dataout<=36'h1fcc9eff0;
			11'h422: dataout<=36'h2f125dc1b;
			11'h423: dataout<=36'h3d9b9c0ca;
			11'h424: dataout<=36'h0fd79fc0f;
			11'h425: dataout<=36'h1f70df04e;
			11'h426: dataout<=36'h2e8e5dcec;
			11'h427: dataout<=36'h3cf5dc234;
			11'h428: dataout<=36'h0fa95fc26;
			11'h429: dataout<=36'h1f165f0aa;
			11'h42a: dataout<=36'h2e0bdddb7;
			11'h42b: dataout<=36'h3c515c396;
			11'h42c: dataout<=36'h0f7b9fc3c;
			11'h42d: dataout<=36'h1ebcdf102;
			11'h42e: dataout<=36'h2d8a9de7b;
			11'h42f: dataout<=36'h3bae1c4f1;
			11'h430: dataout<=36'h0f4e1fc52;
			11'h431: dataout<=36'h1e63df159;
			11'h432: dataout<=36'h2d0a1df3d;
			11'h433: dataout<=36'h3b0c5c643;
			11'h434: dataout<=36'h0f215fc67;
			11'h435: dataout<=36'h1e0c5f1ae;
			11'h436: dataout<=36'h2c8b5dffa;
			11'h437: dataout<=36'h3a6c1c78f;
			11'h438: dataout<=36'h0ef51fc7c;
			11'h439: dataout<=36'h1db59f201;
			11'h43a: dataout<=36'h2c0dde0b3;
			11'h43b: dataout<=36'h39cd1c8d3;
			11'h43c: dataout<=36'h0ec95fc91;
			11'h43d: dataout<=36'h1d601f253;
			11'h43e: dataout<=36'h2b921e169;
			11'h43f: dataout<=36'h392f9ca0f;
			11'h440: dataout<=36'h0e9e1fca5;
			11'h441: dataout<=36'h1d0b1f2a3;
			11'h442: dataout<=36'h2b16de21a;
			11'h443: dataout<=36'h38935cb45;
			11'h444: dataout<=36'h0e735fcb8;
			11'h445: dataout<=36'h1cb75f2ef;
			11'h446: dataout<=36'h2a9d5e2c5;
			11'h447: dataout<=36'h37f89cc74;
			11'h448: dataout<=36'h0e48dfccc;
			11'h449: dataout<=36'h1c641f33d;
			11'h44a: dataout<=36'h2a245e371;
			11'h44b: dataout<=36'h375f1cd9d;
			11'h44c: dataout<=36'h0e1f1fcde;
			11'h44d: dataout<=36'h1c121f386;
			11'h44e: dataout<=36'h29ad1e415;
			11'h44f: dataout<=36'h36c75cebe;
			11'h450: dataout<=36'h0df5dfcf1;
			11'h451: dataout<=36'h1bc11f3d0;
			11'h452: dataout<=36'h29379e4b8;
			11'h453: dataout<=36'h36309cfda;
			11'h454: dataout<=36'h0dccdfd02;
			11'h455: dataout<=36'h1b705f415;
			11'h456: dataout<=36'h28c21e554;
			11'h457: dataout<=36'h359b5d0ef;
			11'h458: dataout<=36'h0da45fd14;
			11'h459: dataout<=36'h1b20df45c;
			11'h45a: dataout<=36'h284e5e5f1;
			11'h45b: dataout<=36'h35079d1fe;
			11'h45c: dataout<=36'h0d7c5fd25;
			11'h45d: dataout<=36'h1ad25f4a0;
			11'h45e: dataout<=36'h27dbde688;
			11'h45f: dataout<=36'h34751d307;
			11'h460: dataout<=36'h0d54dfd35;
			11'h461: dataout<=36'h1a849f4e1;
			11'h462: dataout<=36'h276a5e71a;
			11'h463: dataout<=36'h33e3dd40a;
			11'h464: dataout<=36'h0d2ddfd46;
			11'h465: dataout<=36'h1a37df523;
			11'h466: dataout<=36'h26fa5e7ac;
			11'h467: dataout<=36'h33541d507;
			11'h468: dataout<=36'h0d075fd56;
			11'h469: dataout<=36'h19ec1f562;
			11'h46a: dataout<=36'h268bde839;
			11'h46b: dataout<=36'h32c5dd5ff;
			11'h46c: dataout<=36'h0ce11fd65;
			11'h46d: dataout<=36'h19a09f59f;
			11'h46e: dataout<=36'h261d9e8c1;
			11'h46f: dataout<=36'h32389d6f1;
			11'h470: dataout<=36'h0cbb5fd74;
			11'h471: dataout<=36'h19565f5db;
			11'h472: dataout<=36'h25b0de948;
			11'h473: dataout<=36'h31acdd7de;
			11'h474: dataout<=36'h0c961fd83;
			11'h475: dataout<=36'h190cdf616;
			11'h476: dataout<=36'h25455e9cb;
			11'h477: dataout<=36'h31229d8c6;
			11'h478: dataout<=36'h0c711fd92;
			11'h479: dataout<=36'h18c41f651;
			11'h47a: dataout<=36'h24dadea4e;
			11'h47b: dataout<=36'h30999d9a8;
			11'h47c: dataout<=36'h0c4c9fda0;
			11'h47d: dataout<=36'h187c1f689;
			11'h47e: dataout<=36'h24719eacb;
			11'h47f: dataout<=36'h3011dda86;
			11'h480: dataout<=36'h0c289fdae;
			11'h481: dataout<=36'h18351f6c1;
			11'h482: dataout<=36'h24099eb48;
			11'h483: dataout<=36'h2f8b5db5e;
			11'h484: dataout<=36'h0c04dfdbb;
			11'h485: dataout<=36'h17ee5f6f5;
			11'h486: dataout<=36'h23a1debbe;
			11'h487: dataout<=36'h2f065dc32;
			11'h488: dataout<=36'h0be19fdc8;
			11'h489: dataout<=36'h17a8df72a;
			11'h48a: dataout<=36'h233bdec33;
			11'h48b: dataout<=36'h2e829dd01;
			11'h48c: dataout<=36'h0bbedfdd5;
			11'h48d: dataout<=36'h17645f75d;
			11'h48e: dataout<=36'h22d71eca6;
			11'h48f: dataout<=36'h2dffdddcb;
			11'h490: dataout<=36'h0b9c5fde2;
			11'h491: dataout<=36'h17201f790;
			11'h492: dataout<=36'h22731ed17;
			11'h493: dataout<=36'h2d7edde91;
			11'h494: dataout<=36'h0b7a5fdee;
			11'h495: dataout<=36'h16dd1f7c1;
			11'h496: dataout<=36'h22109ed85;
			11'h497: dataout<=36'h2cfeddf52;
			11'h498: dataout<=36'h0b589fdfa;
			11'h499: dataout<=36'h169a5f7f1;
			11'h49a: dataout<=36'h21ae5edf0;
			11'h49b: dataout<=36'h2c801e00f;
			11'h49c: dataout<=36'h0b375fe06;
			11'h49d: dataout<=36'h16589f820;
			11'h49e: dataout<=36'h214ddee59;
			11'h49f: dataout<=36'h2c02de0c8;
			11'h4a0: dataout<=36'h0b169fe12;
			11'h4a1: dataout<=36'h1617df84f;
			11'h4a2: dataout<=36'h20ee9eec1;
			11'h4a3: dataout<=36'h2b869e17d;
			11'h4a4: dataout<=36'h0af61fe1d;
			11'h4a5: dataout<=36'h15d79f87b;
			11'h4a6: dataout<=36'h208fdef24;
			11'h4a7: dataout<=36'h2b0b9e22d;
			11'h4a8: dataout<=36'h0ad5dfe28;
			11'h4a9: dataout<=36'h1597df8a7;
			11'h4aa: dataout<=36'h20321ef86;
			11'h4ab: dataout<=36'h2a921e2da;
			11'h4ac: dataout<=36'h0ab61fe33;
			11'h4ad: dataout<=36'h1558df8d2;
			11'h4ae: dataout<=36'h1fd55efe7;
			11'h4af: dataout<=36'h2a199e383;
			11'h4b0: dataout<=36'h0a969fe3d;
			11'h4b1: dataout<=36'h151a9f8fb;
			11'h4b2: dataout<=36'h1f799f043;
			11'h4b3: dataout<=36'h29a25e428;
			11'h4b4: dataout<=36'h0a779fe47;
			11'h4b5: dataout<=36'h14dd1f923;
			11'h4b6: dataout<=36'h1f1edf09d;
			11'h4b7: dataout<=36'h292c5e4c9;
			11'h4b8: dataout<=36'h0a58dfe51;
			11'h4b9: dataout<=36'h14a05f94b;
			11'h4ba: dataout<=36'h1ec51f0f7;
			11'h4bb: dataout<=36'h28b79e567;
			11'h4bc: dataout<=36'h0a3a5fe5b;
			11'h4bd: dataout<=36'h1463df973;
			11'h4be: dataout<=36'h1e6c1f14f;
			11'h4bf: dataout<=36'h28441e601;
			11'h4c0: dataout<=36'h0a1c5fe65;
			11'h4c1: dataout<=36'h14289f99a;
			11'h4c2: dataout<=36'h1e149f1a6;
			11'h4c3: dataout<=36'h27d19e698;
			11'h4c4: dataout<=36'h09fedfe6e;
			11'h4c5: dataout<=36'h13ee1f9be;
			11'h4c6: dataout<=36'h1dbe1f1f8;
			11'h4c7: dataout<=36'h27605e72b;
			11'h4c8: dataout<=36'h09e15fe77;
			11'h4c9: dataout<=36'h13b39f9e3;
			11'h4ca: dataout<=36'h1d679f24a;
			11'h4cb: dataout<=36'h26f05e7bb;
			11'h4cc: dataout<=36'h09c45fe80;
			11'h4cd: dataout<=36'h137a1fa06;
			11'h4ce: dataout<=36'h1d129f299;
			11'h4cf: dataout<=36'h26819e848;
			11'h4d0: dataout<=36'h09a7dfe89;
			11'h4d1: dataout<=36'h13419fa2a;
			11'h4d2: dataout<=36'h1cbf5f2e8;
			11'h4d3: dataout<=36'h2613de8d2;
			11'h4d4: dataout<=36'h098b5fe92;
			11'h4d5: dataout<=36'h13091fa4d;
			11'h4d6: dataout<=36'h1c6b9f336;
			11'h4d7: dataout<=36'h25a71e958;
			11'h4d8: dataout<=36'h096f5fe9a;
			11'h4d9: dataout<=36'h12d19fa6d;
			11'h4da: dataout<=36'h1c199f37f;
			11'h4db: dataout<=36'h253bde9dc;
			11'h4dc: dataout<=36'h0953dfea2;
			11'h4dd: dataout<=36'h129b1fa8d;
			11'h4de: dataout<=36'h1bc8df3c7;
			11'h4df: dataout<=36'h24d15ea5c;
			11'h4e0: dataout<=36'h09385feaa;
			11'h4e1: dataout<=36'h12645faad;
			11'h4e2: dataout<=36'h1b77df40e;
			11'h4e3: dataout<=36'h24681eada;
			11'h4e4: dataout<=36'h091d5feb2;
			11'h4e5: dataout<=36'h122edfacd;
			11'h4e6: dataout<=36'h1b289f455;
			11'h4e7: dataout<=36'h24001eb55;
			11'h4e8: dataout<=36'h09029feb9;
			11'h4e9: dataout<=36'h11f9dfaea;
			11'h4ea: dataout<=36'h1ada1f497;
			11'h4eb: dataout<=36'h23991ebcd;
			11'h4ec: dataout<=36'h08e81fec1;
			11'h4ed: dataout<=36'h11c51fb09;
			11'h4ee: dataout<=36'h1a8c1f4db;
			11'h4ef: dataout<=36'h23331ec42;
			11'h4f0: dataout<=36'h08cddfec8;
			11'h4f1: dataout<=36'h11911fb25;
			11'h4f2: dataout<=36'h1a3edf51b;
			11'h4f3: dataout<=36'h22ce5ecb5;
			11'h4f4: dataout<=36'h08b41fecf;
			11'h4f5: dataout<=36'h115ddfb41;
			11'h4f6: dataout<=36'h19f31f55a;
			11'h4f7: dataout<=36'h226a5ed25;
			11'h4f8: dataout<=36'h089a9fed6;
			11'h4f9: dataout<=36'h112b5fb5d;
			11'h4fa: dataout<=36'h19a81f598;
			11'h4fb: dataout<=36'h2207ded92;
			11'h4fc: dataout<=36'h08815fedd;
			11'h4fd: dataout<=36'h10f91fb78;
			11'h4fe: dataout<=36'h195d9f5d5;
			11'h4ff: dataout<=36'h21a61edfd;
			11'h500: dataout<=36'h08685fee3;
			11'h501: dataout<=36'h10c75fb92;
			11'h502: dataout<=36'h1913df60f;
			11'h503: dataout<=36'h21455ee66;
			11'h504: dataout<=36'h084f9feea;
			11'h505: dataout<=36'h10961fbad;
			11'h506: dataout<=36'h18cadf64b;
			11'h507: dataout<=36'h20e5deecc;
			11'h508: dataout<=36'h08371fef0;
			11'h509: dataout<=36'h10659fbc5;
			11'h50a: dataout<=36'h18829f682;
			11'h50b: dataout<=36'h20875ef31;
			11'h50c: dataout<=36'h081f1fef6;
			11'h50d: dataout<=36'h1035dfbdd;
			11'h50e: dataout<=36'h183bdf6b8;
			11'h50f: dataout<=36'h20299ef92;
			11'h510: dataout<=36'h08071fefc;
			11'h511: dataout<=36'h10061fbf5;
			11'h512: dataout<=36'h17f4df6ee;
			11'h513: dataout<=36'h1fcd1eff2;
			11'h514: dataout<=36'h07ef9ff02;
			11'h515: dataout<=36'h0fd75fc0d;
			11'h516: dataout<=36'h17af9f724;
			11'h517: dataout<=36'h1f719f04f;
			11'h518: dataout<=36'h07d85ff08;
			11'h519: dataout<=36'h0fa91fc25;
			11'h51a: dataout<=36'h176adf758;
			11'h51b: dataout<=36'h1f16df0aa;
			11'h51c: dataout<=36'h07c15ff0e;
			11'h51d: dataout<=36'h0f7b5fc3c;
			11'h51e: dataout<=36'h1726df78c;
			11'h51f: dataout<=36'h1ebd5f104;
			11'h520: dataout<=36'h07aa9ff13;
			11'h521: dataout<=36'h0f4e1fc51;
			11'h522: dataout<=36'h16e39f7bb;
			11'h523: dataout<=36'h1e649f15b;
			11'h524: dataout<=36'h0793dff19;
			11'h525: dataout<=36'h0f20dfc68;
			11'h526: dataout<=36'h16a05f7ee;
			11'h527: dataout<=36'h1e0d1f1b0;
			11'h528: dataout<=36'h077d9ff1e;
			11'h529: dataout<=36'h0ef49fc7c;
			11'h52a: dataout<=36'h165e9f81c;
			11'h52b: dataout<=36'h1db65f203;
			11'h52c: dataout<=36'h07679ff23;
			11'h52d: dataout<=36'h0ec8dfc90;
			11'h52e: dataout<=36'h161d5f849;
			11'h52f: dataout<=36'h1d609f255;
			11'h530: dataout<=36'h0751dff28;
			11'h531: dataout<=36'h0e9d9fca4;
			11'h532: dataout<=36'h15dd1f876;
			11'h533: dataout<=36'h1d0b9f2a4;
			11'h534: dataout<=36'h073c5ff2d;
			11'h535: dataout<=36'h0e72dfcb8;
			11'h536: dataout<=36'h159d5f8a2;
			11'h537: dataout<=36'h1cb79f2f2;
			11'h538: dataout<=36'h07271ff32;
			11'h539: dataout<=36'h0e489fccc;
			11'h53a: dataout<=36'h155e9f8ce;
			11'h53b: dataout<=36'h1c649f33e;
			11'h53c: dataout<=36'h07121ff36;
			11'h53d: dataout<=36'h0e1e9fcdd;
			11'h53e: dataout<=36'h15201f8f6;
			11'h53f: dataout<=36'h1c129f388;
			11'h540: dataout<=36'h06fd5ff3b;
			11'h541: dataout<=36'h0df55fcf0;
			11'h542: dataout<=36'h14e29f920;
			11'h543: dataout<=36'h1bc15f3d1;
			11'h544: dataout<=36'h06e8dff3f;
			11'h545: dataout<=36'h0dcc9fd01;
			11'h546: dataout<=36'h14a5df947;
			11'h547: dataout<=36'h1b711f418;
			11'h548: dataout<=36'h06d49ff44;
			11'h549: dataout<=36'h0da41fd14;
			11'h54a: dataout<=36'h1469df970;
			11'h54b: dataout<=36'h1b219f45d;
			11'h54c: dataout<=36'h06c09ff48;
			11'h54d: dataout<=36'h0d7c5fd24;
			11'h54e: dataout<=36'h142e9f995;
			11'h54f: dataout<=36'h1ad31f4a1;
			11'h550: dataout<=36'h06ac9ff4c;
			11'h551: dataout<=36'h0d549fd34;
			11'h552: dataout<=36'h13f35f9ba;
			11'h553: dataout<=36'h1a855f4e3;
			11'h554: dataout<=36'h06991ff50;
			11'h555: dataout<=36'h0d2d9fd44;
			11'h556: dataout<=36'h13b91f9de;
			11'h557: dataout<=36'h1a385f524;
			11'h558: dataout<=36'h06859ff54;
			11'h559: dataout<=36'h0d06dfd54;
			11'h55a: dataout<=36'h137f5fa02;
			11'h55b: dataout<=36'h19ec5f563;
			11'h55c: dataout<=36'h06729ff58;
			11'h55d: dataout<=36'h0ce11fd64;
			11'h55e: dataout<=36'h13471fa25;
			11'h55f: dataout<=36'h19a11f5a1;
			11'h560: dataout<=36'h065f9ff5c;
			11'h561: dataout<=36'h0cbb1fd74;
			11'h562: dataout<=36'h130e9fa48;
			11'h563: dataout<=36'h1956df5de;
			11'h564: dataout<=36'h064cdff60;
			11'h565: dataout<=36'h0c95dfd83;
			11'h566: dataout<=36'h12d71fa6a;
			11'h567: dataout<=36'h190d5f619;
			11'h568: dataout<=36'h063a5ff63;
			11'h569: dataout<=36'h0c70dfd90;
			11'h56a: dataout<=36'h129fdfa88;
			11'h56b: dataout<=36'h18c49f652;
			11'h56c: dataout<=36'h06281ff67;
			11'h56d: dataout<=36'h0c4c9fd9f;
			11'h56e: dataout<=36'h1269dfaa9;
			11'h56f: dataout<=36'h187c9f68b;
			11'h570: dataout<=36'h0615dff6a;
			11'h571: dataout<=36'h0c281fdac;
			11'h572: dataout<=36'h12335fac7;
			11'h573: dataout<=36'h18359f6c2;
			11'h574: dataout<=36'h06041ff6e;
			11'h575: dataout<=36'h0c04dfdbb;
			11'h576: dataout<=36'h11fedfae8;
			11'h577: dataout<=36'h17ef1f6f8;
			11'h578: dataout<=36'h05f25ff71;
			11'h579: dataout<=36'h0be15fdc8;
			11'h57a: dataout<=36'h11c9dfb05;
			11'h57b: dataout<=36'h17a99f72c;
			11'h57c: dataout<=36'h05e0dff74;
			11'h57d: dataout<=36'h0bbe9fdd4;
			11'h57e: dataout<=36'h1195dfb21;
			11'h57f: dataout<=36'h1764df760;
			11'h580: dataout<=36'h05cf9ff77;
			11'h581: dataout<=36'h0b9c1fde0;
			11'h582: dataout<=36'h11625fb3c;
			11'h583: dataout<=36'h1720df792;
			11'h584: dataout<=36'h05be9ff7a;
			11'h585: dataout<=36'h0b7a5fded;
			11'h586: dataout<=36'h11301fb59;
			11'h587: dataout<=36'h16dd9f7c3;
			11'h588: dataout<=36'h05ad9ff7d;
			11'h589: dataout<=36'h0b585fdf9;
			11'h58a: dataout<=36'h10fd5fb74;
			11'h58b: dataout<=36'h169b1f7f3;
			11'h58c: dataout<=36'h059cdff80;
			11'h58d: dataout<=36'h0b36dfe05;
			11'h58e: dataout<=36'h10cb5fb8e;
			11'h58f: dataout<=36'h16595f822;
			11'h590: dataout<=36'h058c5ff83;
			11'h591: dataout<=36'h0b161fe10;
			11'h592: dataout<=36'h109a5fba8;
			11'h593: dataout<=36'h16181f850;
			11'h594: dataout<=36'h057c1ff86;
			11'h595: dataout<=36'h0af59fe1c;
			11'h596: dataout<=36'h1069dfbc2;
			11'h597: dataout<=36'h15d7df87d;
			11'h598: dataout<=36'h056c1ff89;
			11'h599: dataout<=36'h0ad59fe27;
			11'h59a: dataout<=36'h103a1fbdb;
			11'h59b: dataout<=36'h15985f8a9;
			11'h59c: dataout<=36'h055c1ff8b;
			11'h59d: dataout<=36'h0ab5dfe31;
			11'h59e: dataout<=36'h100a9fbf2;
			11'h59f: dataout<=36'h15595f8d3;
			11'h5a0: dataout<=36'h054c5ff8e;
			11'h5a1: dataout<=36'h0a965fe3c;
			11'h5a2: dataout<=36'h0fdb9fc0a;
			11'h5a3: dataout<=36'h151b1f8fd;
			11'h5a4: dataout<=36'h053cdff91;
			11'h5a5: dataout<=36'h0a775fe47;
			11'h5a6: dataout<=36'h0fad5fc22;
			11'h5a7: dataout<=36'h14dd9f926;
			11'h5a8: dataout<=36'h052d5ff93;
			11'h5a9: dataout<=36'h0a589fe50;
			11'h5aa: dataout<=36'h0f7f5fc37;
			11'h5ab: dataout<=36'h14a0df94e;
			11'h5ac: dataout<=36'h051e1ff96;
			11'h5ad: dataout<=36'h0a3a1fe5b;
			11'h5ae: dataout<=36'h0f51dfc4f;
			11'h5af: dataout<=36'h14649f975;
			11'h5b0: dataout<=36'h050f1ff98;
			11'h5b1: dataout<=36'h0a1c1fe64;
			11'h5b2: dataout<=36'h0f251fc64;
			11'h5b3: dataout<=36'h14295f99b;
			11'h5b4: dataout<=36'h05005ff9a;
			11'h5b5: dataout<=36'h09fedfe6c;
			11'h5b6: dataout<=36'h0ef95fc77;
			11'h5b7: dataout<=36'h13ee5f9c1;
			11'h5b8: dataout<=36'h04f19ff9d;
			11'h5b9: dataout<=36'h09e15fe77;
			11'h5ba: dataout<=36'h0ecd5fc8e;
			11'h5bb: dataout<=36'h13b45f9e5;
			11'h5bc: dataout<=36'h04e31ff9f;
			11'h5bd: dataout<=36'h09c45fe7f;
			11'h5be: dataout<=36'h0ea1dfca1;
			11'h5bf: dataout<=36'h137adfa09;
			11'h5c0: dataout<=36'h04d49ffa1;
			11'h5c1: dataout<=36'h09a75fe88;
			11'h5c2: dataout<=36'h0e769fcb5;
			11'h5c3: dataout<=36'h13421fa2c;
			11'h5c4: dataout<=36'h04c65ffa3;
			11'h5c5: dataout<=36'h098b1fe90;
			11'h5c6: dataout<=36'h0e4c5fcc7;
			11'h5c7: dataout<=36'h1309dfa4e;
			11'h5c8: dataout<=36'h04b85ffa5;
			11'h5c9: dataout<=36'h096f1fe98;
			11'h5ca: dataout<=36'h0e229fcd9;
			11'h5cb: dataout<=36'h12d25fa6f;
			11'h5cc: dataout<=36'h04aa9ffa7;
			11'h5cd: dataout<=36'h09539fea0;
			11'h5ce: dataout<=36'h0df95fcec;
			11'h5cf: dataout<=36'h129b5fa8f;
			11'h5d0: dataout<=36'h049cdffa9;
			11'h5d1: dataout<=36'h09381fea8;
			11'h5d2: dataout<=36'h0dd05fcfd;
			11'h5d3: dataout<=36'h1264dfaaf;
			11'h5d4: dataout<=36'h048f5ffab;
			11'h5d5: dataout<=36'h091d1feb0;
			11'h5d6: dataout<=36'h0da81fd0f;
			11'h5d7: dataout<=36'h122f5face;
			11'h5d8: dataout<=36'h0481dffad;
			11'h5d9: dataout<=36'h09025feb8;
			11'h5da: dataout<=36'h0d7fdfd21;
			11'h5db: dataout<=36'h11fa1faec;
			11'h5dc: dataout<=36'h04749ffaf;
			11'h5dd: dataout<=36'h08e7dfec0;
			11'h5de: dataout<=36'h0d585fd32;
			11'h5df: dataout<=36'h11c59fb0a;
			11'h5e0: dataout<=36'h04679ffb1;
			11'h5e1: dataout<=36'h08cddfec7;
			11'h5e2: dataout<=36'h0d315fd42;
			11'h5e3: dataout<=36'h11919fb27;
			11'h5e4: dataout<=36'h045a9ffb3;
			11'h5e5: dataout<=36'h08b3dfecf;
			11'h5e6: dataout<=36'h0d0a9fd54;
			11'h5e7: dataout<=36'h115e5fb43;
			11'h5e8: dataout<=36'h044ddffb4;
			11'h5e9: dataout<=36'h089a5fed4;
			11'h5ea: dataout<=36'h0ce45fd60;
			11'h5eb: dataout<=36'h112b9fb5f;
			11'h5ec: dataout<=36'h04411ffb6;
			11'h5ed: dataout<=36'h08811fedc;
			11'h5ee: dataout<=36'h0cbe9fd71;
			11'h5ef: dataout<=36'h10f95fb7a;
			11'h5f0: dataout<=36'h04349ffb8;
			11'h5f1: dataout<=36'h08681fee3;
			11'h5f2: dataout<=36'h0c991fd81;
			11'h5f3: dataout<=36'h10c7dfb94;
			11'h5f4: dataout<=36'h04281ffb9;
			11'h5f5: dataout<=36'h084f1fee8;
			11'h5f6: dataout<=36'h0c73dfd8d;
			11'h5f7: dataout<=36'h10969fbae;
			11'h5f8: dataout<=36'h041c1ffbb;
			11'h5f9: dataout<=36'h08371feef;
			11'h5fa: dataout<=36'h0c4fdfd9d;
			11'h5fb: dataout<=36'h10661fbc7;
			11'h5fc: dataout<=36'h040fdffbc;
			11'h5fd: dataout<=36'h081e9fef5;
			11'h5fe: dataout<=36'h0c2b5fdaa;
			11'h5ff: dataout<=36'h10365fbe0;
			11'h600: dataout<=36'h0403dffbe;
			11'h601: dataout<=36'h08069fefc;
			11'h602: dataout<=36'h0c075fdb9;
			11'h603: dataout<=36'h1006dfbf8;
			11'h604: dataout<=36'h03f81ffbf;
			11'h605: dataout<=36'h07ef1ff00;
			11'h606: dataout<=36'h0be45fdc4;
			11'h607: dataout<=36'h0fd7dfc10;
			11'h608: dataout<=36'h03ec9ffc1;
			11'h609: dataout<=36'h07d85ff07;
			11'h60a: dataout<=36'h0bc21fdd2;
			11'h60b: dataout<=36'h0fa99fc27;
			11'h60c: dataout<=36'h03e0dffc2;
			11'h60d: dataout<=36'h07c0dff0c;
			11'h60e: dataout<=36'h0b9edfdde;
			11'h60f: dataout<=36'h0f7bdfc3d;
			11'h610: dataout<=36'h03d59ffc4;
			11'h611: dataout<=36'h07aa5ff13;
			11'h612: dataout<=36'h0b7d5fdec;
			11'h613: dataout<=36'h0f4e5fc53;
			11'h614: dataout<=36'h03ca5ffc5;
			11'h615: dataout<=36'h0793dff18;
			11'h616: dataout<=36'h0b5b9fdf8;
			11'h617: dataout<=36'h0f219fc68;
			11'h618: dataout<=36'h03bf1ffc6;
			11'h619: dataout<=36'h077d5ff1c;
			11'h61a: dataout<=36'h0b39dfe02;
			11'h61b: dataout<=36'h0ef55fc7d;
			11'h61c: dataout<=36'h03b41ffc8;
			11'h61d: dataout<=36'h07675ff23;
			11'h61e: dataout<=36'h0b191fe10;
			11'h61f: dataout<=36'h0ec99fc92;
			11'h620: dataout<=36'h03a91ffc9;
			11'h621: dataout<=36'h07515ff27;
			11'h622: dataout<=36'h0af81fe1a;
			11'h623: dataout<=36'h0e9e5fca6;
			11'h624: dataout<=36'h039e5ffca;
			11'h625: dataout<=36'h073bdff2c;
			11'h626: dataout<=36'h0ad81fe25;
			11'h627: dataout<=36'h0e739fcb9;
			11'h628: dataout<=36'h0393dffcb;
			11'h629: dataout<=36'h07271ff30;
			11'h62a: dataout<=36'h0ab8dfe2f;
			11'h62b: dataout<=36'h0e491fccd;
			11'h62c: dataout<=36'h03895ffcc;
			11'h62d: dataout<=36'h07121ff34;
			11'h62e: dataout<=36'h0a995fe39;
			11'h62f: dataout<=36'h0e1f5fcdf;
			11'h630: dataout<=36'h037edffce;
			11'h631: dataout<=36'h06fd1ff3b;
			11'h632: dataout<=36'h0a79dfe46;
			11'h633: dataout<=36'h0df61fcf2;
			11'h634: dataout<=36'h03749ffcf;
			11'h635: dataout<=36'h06e89ff3f;
			11'h636: dataout<=36'h0a5b5fe50;
			11'h637: dataout<=36'h0dcd1fd03;
			11'h638: dataout<=36'h036a5ffd0;
			11'h639: dataout<=36'h06d41ff43;
			11'h63a: dataout<=36'h0a3c9fe59;
			11'h63b: dataout<=36'h0da49fd15;
			11'h63c: dataout<=36'h03605ffd1;
			11'h63d: dataout<=36'h06c01ff47;
			11'h63e: dataout<=36'h0a1e9fe62;
			11'h63f: dataout<=36'h0d7c9fd26;
			11'h640: dataout<=36'h03569ffd2;
			11'h641: dataout<=36'h06ac9ff4b;
			11'h642: dataout<=36'h0a015fe6b;
			11'h643: dataout<=36'h0d551fd36;
			11'h644: dataout<=36'h034c9ffd3;
			11'h645: dataout<=36'h06989ff4f;
			11'h646: dataout<=36'h09e39fe74;
			11'h647: dataout<=36'h0d2e1fd47;
			11'h648: dataout<=36'h0342dffd4;
			11'h649: dataout<=36'h06851ff53;
			11'h64a: dataout<=36'h09c65fe7d;
			11'h64b: dataout<=36'h0d079fd57;
			11'h64c: dataout<=36'h03395ffd5;
			11'h64d: dataout<=36'h06721ff57;
			11'h64e: dataout<=36'h09a9dfe86;
			11'h64f: dataout<=36'h0ce15fd66;
			11'h650: dataout<=36'h032fdffd6;
			11'h651: dataout<=36'h065f1ff5b;
			11'h652: dataout<=36'h098d5fe8f;
			11'h653: dataout<=36'h0cbb9fd75;
			11'h654: dataout<=36'h03269ffd7;
			11'h655: dataout<=36'h064cdff5f;
			11'h656: dataout<=36'h09721fe98;
			11'h657: dataout<=36'h0c965fd84;
			11'h658: dataout<=36'h031d5ffd8;
			11'h659: dataout<=36'h063a5ff63;
			11'h65a: dataout<=36'h09565fea0;
			11'h65b: dataout<=36'h0c715fd93;
			11'h65c: dataout<=36'h03141ffd9;
			11'h65d: dataout<=36'h0627dff67;
			11'h65e: dataout<=36'h093a9fea9;
			11'h65f: dataout<=36'h0c4cdfda1;
			11'h660: dataout<=36'h030b1ffd9;
			11'h661: dataout<=36'h0615dff68;
			11'h662: dataout<=36'h091f9fead;
			11'h663: dataout<=36'h0c28dfdaf;
			11'h664: dataout<=36'h03021ffda;
			11'h665: dataout<=36'h0603dff6c;
			11'h666: dataout<=36'h09049feb6;
			11'h667: dataout<=36'h0c051fdbc;
			11'h668: dataout<=36'h02f95ffdb;
			11'h669: dataout<=36'h05f25ff70;
			11'h66a: dataout<=36'h08ea5febe;
			11'h66b: dataout<=36'h0be1dfdc9;
			11'h66c: dataout<=36'h02f09ffdc;
			11'h66d: dataout<=36'h05e0dff73;
			11'h66e: dataout<=36'h08d05fec5;
			11'h66f: dataout<=36'h0bbf1fdd6;
			11'h670: dataout<=36'h02e7dffdd;
			11'h671: dataout<=36'h05cf5ff77;
			11'h672: dataout<=36'h08b61fecd;
			11'h673: dataout<=36'h0b9c9fde3;
			11'h674: dataout<=36'h02df5ffdd;
			11'h675: dataout<=36'h05be5ff78;
			11'h676: dataout<=36'h089c9fed2;
			11'h677: dataout<=36'h0b7a9fdef;
			11'h678: dataout<=36'h02d6dffde;
			11'h679: dataout<=36'h05ad5ff7c;
			11'h67a: dataout<=36'h08831feda;
			11'h67b: dataout<=36'h0b58dfdfb;
			11'h67c: dataout<=36'h02ce9ffdf;
			11'h67d: dataout<=36'h059cdff7f;
			11'h67e: dataout<=36'h086a5fee0;
			11'h67f: dataout<=36'h0b379fe07;
			11'h680: dataout<=36'h02c65ffe0;
			11'h681: dataout<=36'h058c5ff83;
			11'h682: dataout<=36'h08519fee8;
			11'h683: dataout<=36'h0b16dfe13;
			11'h684: dataout<=36'h02be1ffe0;
			11'h685: dataout<=36'h057bdff84;
			11'h686: dataout<=36'h08391feec;
			11'h687: dataout<=36'h0af65fe1e;
			11'h688: dataout<=36'h02b61ffe1;
			11'h689: dataout<=36'h056bdff88;
			11'h68a: dataout<=36'h08211fef4;
			11'h68b: dataout<=36'h0ad61fe29;
			11'h68c: dataout<=36'h02ae1ffe2;
			11'h68d: dataout<=36'h055bdff8b;
			11'h68e: dataout<=36'h08091fefb;
			11'h68f: dataout<=36'h0ab65fe34;
			11'h690: dataout<=36'h02a61ffe2;
			11'h691: dataout<=36'h054bdff8c;
			11'h692: dataout<=36'h07f11fefe;
			11'h693: dataout<=36'h0a96dfe3e;
			11'h694: dataout<=36'h029e5ffe3;
			11'h695: dataout<=36'h053c5ff90;
			11'h696: dataout<=36'h07d9dff06;
			11'h697: dataout<=36'h0a77dfe48;
			11'h698: dataout<=36'h02969ffe4;
			11'h699: dataout<=36'h052cdff93;
			11'h69a: dataout<=36'h07c29ff0c;
			11'h69b: dataout<=36'h0a591fe52;
			11'h69c: dataout<=36'h028f1ffe4;
			11'h69d: dataout<=36'h051ddff94;
			11'h69e: dataout<=36'h07ac1ff10;
			11'h69f: dataout<=36'h0a3a9fe5c;
			11'h6a0: dataout<=36'h02879ffe5;
			11'h6a1: dataout<=36'h050edff97;
			11'h6a2: dataout<=36'h07959ff16;
			11'h6a3: dataout<=36'h0a1c9fe66;
			11'h6a4: dataout<=36'h02801ffe5;
			11'h6a5: dataout<=36'h04ffdff98;
			11'h6a6: dataout<=36'h077f1ff1a;
			11'h6a7: dataout<=36'h09ff1fe6f;
			11'h6a8: dataout<=36'h0278dffe6;
			11'h6a9: dataout<=36'h04f19ff9c;
			11'h6aa: dataout<=36'h0769dff21;
			11'h6ab: dataout<=36'h09e19fe78;
			11'h6ac: dataout<=36'h02719ffe7;
			11'h6ad: dataout<=36'h04e31ff9f;
			11'h6ae: dataout<=36'h07541ff27;
			11'h6af: dataout<=36'h09c49fe81;
			11'h6b0: dataout<=36'h026a5ffe7;
			11'h6b1: dataout<=36'h04d49ffa0;
			11'h6b2: dataout<=36'h073e5ff2a;
			11'h6b3: dataout<=36'h09a81fe8a;
			11'h6b4: dataout<=36'h02631ffe8;
			11'h6b5: dataout<=36'h04c61ffa3;
			11'h6b6: dataout<=36'h07289ff30;
			11'h6b7: dataout<=36'h098b9fe93;
			11'h6b8: dataout<=36'h025c1ffe8;
			11'h6b9: dataout<=36'h04b81ffa4;
			11'h6ba: dataout<=36'h07139ff33;
			11'h6bb: dataout<=36'h096f9fe9b;
			11'h6bc: dataout<=36'h02551ffe9;
			11'h6bd: dataout<=36'h04aa1ffa7;
			11'h6be: dataout<=36'h06fe9ff39;
			11'h6bf: dataout<=36'h09541fea3;
			11'h6c0: dataout<=36'h024e5ffe9;
			11'h6c1: dataout<=36'h049c9ffa8;
			11'h6c2: dataout<=36'h06ea5ff3c;
			11'h6c3: dataout<=36'h09389feab;
			11'h6c4: dataout<=36'h02479ffea;
			11'h6c5: dataout<=36'h048f1ffab;
			11'h6c6: dataout<=36'h06d61ff42;
			11'h6c7: dataout<=36'h091d9feb3;
			11'h6c8: dataout<=36'h0240dffea;
			11'h6c9: dataout<=36'h04819ffac;
			11'h6ca: dataout<=36'h06c1dff45;
			11'h6cb: dataout<=36'h0902dfeba;
			11'h6cc: dataout<=36'h023a5ffeb;
			11'h6cd: dataout<=36'h04749ffaf;
			11'h6ce: dataout<=36'h06ae5ff4b;
			11'h6cf: dataout<=36'h08e85fec2;
			11'h6d0: dataout<=36'h02339ffeb;
			11'h6d1: dataout<=36'h04671ffb0;
			11'h6d2: dataout<=36'h069a1ff4e;
			11'h6d3: dataout<=36'h08ce1fec9;
			11'h6d4: dataout<=36'h022d1ffec;
			11'h6d5: dataout<=36'h045a1ffb3;
			11'h6d6: dataout<=36'h0686dff54;
			11'h6d7: dataout<=36'h08b45fed0;
			11'h6d8: dataout<=36'h0226dffec;
			11'h6d9: dataout<=36'h044d9ffb3;
			11'h6da: dataout<=36'h06741ff55;
			11'h6db: dataout<=36'h089adfed7;
			11'h6dc: dataout<=36'h02209ffec;
			11'h6dd: dataout<=36'h04411ffb4;
			11'h6de: dataout<=36'h06615ff58;
			11'h6df: dataout<=36'h08819fede;
			11'h6e0: dataout<=36'h021a5ffed;
			11'h6e1: dataout<=36'h04349ffb7;
			11'h6e2: dataout<=36'h064e9ff5e;
			11'h6e3: dataout<=36'h08689fee4;
			11'h6e4: dataout<=36'h02141ffed;
			11'h6e5: dataout<=36'h04281ffb8;
			11'h6e6: dataout<=36'h063bdff60;
			11'h6e7: dataout<=36'h084fdfeeb;
			11'h6e8: dataout<=36'h020ddffee;
			11'h6e9: dataout<=36'h041b9ffbb;
			11'h6ea: dataout<=36'h06291ff66;
			11'h6eb: dataout<=36'h08375fef1;
			11'h6ec: dataout<=36'h0207dffee;
			11'h6ed: dataout<=36'h040f9ffbc;
			11'h6ee: dataout<=36'h06171ff69;
			11'h6ef: dataout<=36'h081f5fef7;
			11'h6f0: dataout<=36'h0201dffee;
			11'h6f1: dataout<=36'h04039ffbc;
			11'h6f2: dataout<=36'h06051ff6a;
			11'h6f3: dataout<=36'h08075fefd;
			11'h6f4: dataout<=36'h01fc1ffef;
			11'h6f5: dataout<=36'h03f81ffbf;
			11'h6f6: dataout<=36'h05f3dff6f;
			11'h6f7: dataout<=36'h07efdff03;
			11'h6f8: dataout<=36'h01f61ffef;
			11'h6f9: dataout<=36'h03ec1ffc0;
			11'h6fa: dataout<=36'h05e1dff72;
			11'h6fb: dataout<=36'h07d89ff09;
			11'h6fc: dataout<=36'h01f05ffef;
			11'h6fd: dataout<=36'h03e09ffc0;
			11'h6fe: dataout<=36'h05d09ff73;
			11'h6ff: dataout<=36'h07c19ff0f;
			11'h700: dataout<=36'h01ea9fff0;
			11'h701: dataout<=36'h03d51ffc3;
			11'h702: dataout<=36'h05bf5ff79;
			11'h703: dataout<=36'h07aadff14;
			11'h704: dataout<=36'h01e51fff0;
			11'h705: dataout<=36'h03ca1ffc4;
			11'h706: dataout<=36'h05aedff7b;
			11'h707: dataout<=36'h07941ff1a;
			11'h708: dataout<=36'h01df9fff0;
			11'h709: dataout<=36'h03bf1ffc4;
			11'h70a: dataout<=36'h059e5ff7c;
			11'h70b: dataout<=36'h077ddff1f;
			11'h70c: dataout<=36'h01d9dfff1;
			11'h70d: dataout<=36'h03b39ffc7;
			11'h70e: dataout<=36'h058d1ff82;
			11'h70f: dataout<=36'h0767dff24;
			11'h710: dataout<=36'h01d49fff1;
			11'h711: dataout<=36'h03a91ffc8;
			11'h712: dataout<=36'h057d5ff84;
			11'h713: dataout<=36'h07521ff29;
			11'h714: dataout<=36'h01cf1fff1;
			11'h715: dataout<=36'h039e1ffc8;
			11'h716: dataout<=36'h056cdff85;
			11'h717: dataout<=36'h073c9ff2e;
			11'h718: dataout<=36'h01c9dfff2;
			11'h719: dataout<=36'h03939ffcb;
			11'h71a: dataout<=36'h055d1ff8a;
			11'h71b: dataout<=36'h07275ff33;
			11'h71c: dataout<=36'h01c49fff2;
			11'h71d: dataout<=36'h03891ffcb;
			11'h71e: dataout<=36'h054d5ff8b;
			11'h71f: dataout<=36'h07125ff37;
			11'h720: dataout<=36'h01bf5fff2;
			11'h721: dataout<=36'h037e9ffcc;
			11'h722: dataout<=36'h053d9ff8e;
			11'h723: dataout<=36'h06fd9ff3c;
			11'h724: dataout<=36'h01ba1fff3;
			11'h725: dataout<=36'h03741ffcf;
			11'h726: dataout<=36'h052e1ff93;
			11'h727: dataout<=36'h06e91ff40;
			11'h728: dataout<=36'h01b51fff3;
			11'h729: dataout<=36'h036a1ffcf;
			11'h72a: dataout<=36'h051f1ff94;
			11'h72b: dataout<=36'h06d4dff45;
			11'h72c: dataout<=36'h01b01fff3;
			11'h72d: dataout<=36'h03601ffd0;
			11'h72e: dataout<=36'h05101ff96;
			11'h72f: dataout<=36'h06c0dff49;
			11'h730: dataout<=36'h01ab1fff3;
			11'h731: dataout<=36'h03561ffd0;
			11'h732: dataout<=36'h05011ff97;
			11'h733: dataout<=36'h06acdff4d;
			11'h734: dataout<=36'h01a65fff4;
			11'h735: dataout<=36'h034c9ffd3;
			11'h736: dataout<=36'h04f2dff9c;
			11'h737: dataout<=36'h06995ff51;
			11'h738: dataout<=36'h01a15fff4;
			11'h739: dataout<=36'h03429ffd3;
			11'h73a: dataout<=36'h04e3dff9d;
			11'h73b: dataout<=36'h0685dff55;
			11'h73c: dataout<=36'h019c9fff4;
			11'h73d: dataout<=36'h03391ffd4;
			11'h73e: dataout<=36'h04d59ff9f;
			11'h73f: dataout<=36'h0672dff59;
			11'h740: dataout<=36'h0197dfff4;
			11'h741: dataout<=36'h032f9ffd4;
			11'h742: dataout<=36'h04c75ffa0;
			11'h743: dataout<=36'h065fdff5d;
			11'h744: dataout<=36'h01931fff5;
			11'h745: dataout<=36'h03261ffd7;
			11'h746: dataout<=36'h04b91ffa5;
			11'h747: dataout<=36'h064d1ff61;
			11'h748: dataout<=36'h018e9fff5;
			11'h749: dataout<=36'h031d1ffd7;
			11'h74a: dataout<=36'h04ab9ffa6;
			11'h74b: dataout<=36'h063a9ff64;
			11'h74c: dataout<=36'h0189dfff5;
			11'h74d: dataout<=36'h03139ffd8;
			11'h74e: dataout<=36'h049d5ffa8;
			11'h74f: dataout<=36'h06285ff68;
			11'h750: dataout<=36'h01855fff5;
			11'h751: dataout<=36'h030a9ffd8;
			11'h752: dataout<=36'h048fdffa8;
			11'h753: dataout<=36'h06161ff6b;
			11'h754: dataout<=36'h0180dfff5;
			11'h755: dataout<=36'h03019ffd8;
			11'h756: dataout<=36'h04825ffa9;
			11'h757: dataout<=36'h06045ff6f;
			11'h758: dataout<=36'h017c9fff6;
			11'h759: dataout<=36'h02f91ffdb;
			11'h75a: dataout<=36'h04759ffae;
			11'h75b: dataout<=36'h05f29ff72;
			11'h75c: dataout<=36'h01781fff6;
			11'h75d: dataout<=36'h02f01ffdb;
			11'h75e: dataout<=36'h04681ffaf;
			11'h75f: dataout<=36'h05e11ff75;
			11'h760: dataout<=36'h0173dfff6;
			11'h761: dataout<=36'h02e79ffdc;
			11'h762: dataout<=36'h045b5ffb1;
			11'h763: dataout<=36'h05cfdff78;
			11'h764: dataout<=36'h016f9fff6;
			11'h765: dataout<=36'h02df1ffdc;
			11'h766: dataout<=36'h044e9ffb2;
			11'h767: dataout<=36'h05bedff7b;
			11'h768: dataout<=36'h016b5fff6;
			11'h769: dataout<=36'h02d69ffdc;
			11'h76a: dataout<=36'h0441dffb2;
			11'h76b: dataout<=36'h05addff7e;
			11'h76c: dataout<=36'h01671fff7;
			11'h76d: dataout<=36'h02ce1ffdf;
			11'h76e: dataout<=36'h04351ffb7;
			11'h76f: dataout<=36'h059d1ff81;
			11'h770: dataout<=36'h01631fff7;
			11'h771: dataout<=36'h02c61ffdf;
			11'h772: dataout<=36'h04291ffb8;
			11'h773: dataout<=36'h058c9ff84;
			11'h774: dataout<=36'h015edfff7;
			11'h775: dataout<=36'h02bd9ffdf;
			11'h776: dataout<=36'h041c5ffb8;
			11'h777: dataout<=36'h057c5ff87;
			11'h778: dataout<=36'h015adfff7;
			11'h779: dataout<=36'h02b59ffe0;
			11'h77a: dataout<=36'h04105ffba;
			11'h77b: dataout<=36'h056c5ff8a;
			11'h77c: dataout<=36'h0156dfff7;
			11'h77d: dataout<=36'h02ad9ffe0;
			11'h77e: dataout<=36'h04045ffbb;
			11'h77f: dataout<=36'h055c5ff8c;
			11'h780: dataout<=36'h000000000;
			11'h781: dataout<=36'h000000000;
			11'h782: dataout<=36'h000000000;
			11'h783: dataout<=36'h000000000;
			11'h784: dataout<=36'h000000000;
			11'h785: dataout<=36'h000000000;
			11'h786: dataout<=36'h000000000;
			11'h787: dataout<=36'h000000000;
			11'h788: dataout<=36'h000000000;
			11'h789: dataout<=36'h000000000;
			11'h78a: dataout<=36'h000000000;
			11'h78b: dataout<=36'h000000000;
			11'h78c: dataout<=36'h000000000;
			11'h78d: dataout<=36'h000000000;
			11'h78e: dataout<=36'h000000000;
			11'h78f: dataout<=36'h000000000;
			11'h790: dataout<=36'h000000000;
			11'h791: dataout<=36'h000000000;
			11'h792: dataout<=36'h000000000;
			11'h793: dataout<=36'h000000000;
			11'h794: dataout<=36'h000000000;
			11'h795: dataout<=36'h000000000;
			11'h796: dataout<=36'h000000000;
			11'h797: dataout<=36'h000000000;
			11'h798: dataout<=36'h000000000;
			11'h799: dataout<=36'h000000000;
			11'h79a: dataout<=36'h000000000;
			11'h79b: dataout<=36'h000000000;
			11'h79c: dataout<=36'h000000000;
			11'h79d: dataout<=36'h000000000;
			11'h79e: dataout<=36'h000000000;
			11'h79f: dataout<=36'h000000000;
			11'h7a0: dataout<=36'h000000000;
			11'h7a1: dataout<=36'h000000000;
			11'h7a2: dataout<=36'h000000000;
			11'h7a3: dataout<=36'h000000000;
			11'h7a4: dataout<=36'h000000000;
			11'h7a5: dataout<=36'h000000000;
			11'h7a6: dataout<=36'h000000000;
			11'h7a7: dataout<=36'h000000000;
			11'h7a8: dataout<=36'h000000000;
			11'h7a9: dataout<=36'h000000000;
			11'h7aa: dataout<=36'h000000000;
			11'h7ab: dataout<=36'h000000000;
			11'h7ac: dataout<=36'h000000000;
			11'h7ad: dataout<=36'h000000000;
			11'h7ae: dataout<=36'h000000000;
			11'h7af: dataout<=36'h000000000;
			11'h7b0: dataout<=36'h000000000;
			11'h7b1: dataout<=36'h000000000;
			11'h7b2: dataout<=36'h000000000;
			11'h7b3: dataout<=36'h000000000;
			11'h7b4: dataout<=36'h000000000;
			11'h7b5: dataout<=36'h000000000;
			11'h7b6: dataout<=36'h000000000;
			11'h7b7: dataout<=36'h000000000;
			11'h7b8: dataout<=36'h000000000;
			11'h7b9: dataout<=36'h000000000;
			11'h7ba: dataout<=36'h000000000;
			11'h7bb: dataout<=36'h000000000;
			11'h7bc: dataout<=36'h000000000;
			11'h7bd: dataout<=36'h000000000;
			11'h7be: dataout<=36'h000000000;
			11'h7bf: dataout<=36'h000000000;
			11'h7c0: dataout<=36'h000000000;
			11'h7c1: dataout<=36'h000000000;
			11'h7c2: dataout<=36'h000000000;
			11'h7c3: dataout<=36'h000000000;
			11'h7c4: dataout<=36'h000000000;
			11'h7c5: dataout<=36'h000000000;
			11'h7c6: dataout<=36'h000000000;
			11'h7c7: dataout<=36'h000000000;
			11'h7c8: dataout<=36'h000000000;
			11'h7c9: dataout<=36'h000000000;
			11'h7ca: dataout<=36'h000000000;
			11'h7cb: dataout<=36'h000000000;
			11'h7cc: dataout<=36'h000000000;
			11'h7cd: dataout<=36'h000000000;
			11'h7ce: dataout<=36'h000000000;
			11'h7cf: dataout<=36'h000000000;
			11'h7d0: dataout<=36'h000000000;
			11'h7d1: dataout<=36'h000000000;
			11'h7d2: dataout<=36'h000000000;
			11'h7d3: dataout<=36'h000000000;
			11'h7d4: dataout<=36'h000000000;
			11'h7d5: dataout<=36'h000000000;
			11'h7d6: dataout<=36'h000000000;
			11'h7d7: dataout<=36'h000000000;
			11'h7d8: dataout<=36'h000000000;
			11'h7d9: dataout<=36'h000000000;
			11'h7da: dataout<=36'h000000000;
			11'h7db: dataout<=36'h000000000;
			11'h7dc: dataout<=36'h000000000;
			11'h7dd: dataout<=36'h000000000;
			11'h7de: dataout<=36'h000000000;
			11'h7df: dataout<=36'h000000000;
			11'h7e0: dataout<=36'h000000000;
			11'h7e1: dataout<=36'h000000000;
			11'h7e2: dataout<=36'h000000000;
			11'h7e3: dataout<=36'h000000000;
			11'h7e4: dataout<=36'h000000000;
			11'h7e5: dataout<=36'h000000000;
			11'h7e6: dataout<=36'h000000000;
			11'h7e7: dataout<=36'h000000000;
			11'h7e8: dataout<=36'h000000000;
			11'h7e9: dataout<=36'h000000000;
			11'h7ea: dataout<=36'h000000000;
			11'h7eb: dataout<=36'h000000000;
			11'h7ec: dataout<=36'h000000000;
			11'h7ed: dataout<=36'h000000000;
			11'h7ee: dataout<=36'h000000000;
			11'h7ef: dataout<=36'h000000000;
			11'h7f0: dataout<=36'h000000000;
			11'h7f1: dataout<=36'h000000000;
			11'h7f2: dataout<=36'h000000000;
			11'h7f3: dataout<=36'h000000000;
			11'h7f4: dataout<=36'h000000000;
			11'h7f5: dataout<=36'h000000000;
			11'h7f6: dataout<=36'h000000000;
			11'h7f7: dataout<=36'h000000000;
			11'h7f8: dataout<=36'h000000000;
			11'h7f9: dataout<=36'h000000000;
			11'h7fa: dataout<=36'h000000000;
			11'h7fb: dataout<=36'h000000000;
			11'h7fc: dataout<=36'h000000000;
			11'h7fd: dataout<=36'h000000000;
			11'h7fe: dataout<=36'h000000000;
			11'h7ff: dataout<=36'h000000000;
		endcase
	end
endmodule

