module nco_rom_4ch_fc2400_fs5859 (clock,addr,dataout);
	input clock;
	input [10:0] addr;
	output reg signed [35:0] dataout;
	always @(posedge clock) begin
		case (addr)
			11'h000: dataout<=36'h460265360;
			11'h001: dataout<=36'h8ac84cda9;
			11'h002: dataout<=36'h7e4045447;
			11'h003: dataout<=36'ha1d4ea538;
			11'h004: dataout<=36'h4694a54e0;
			11'h005: dataout<=36'h8a3d4c8a4;
			11'h006: dataout<=36'h7de5c5c5c;
			11'h007: dataout<=36'ha3b469d41;
			11'h008: dataout<=36'h472665664;
			11'h009: dataout<=36'h89b5cc399;
			11'h00a: dataout<=36'h7d830646a;
			11'h00b: dataout<=36'ha59ea9574;
			11'h00c: dataout<=36'h47b7657ea;
			11'h00d: dataout<=36'h89320be8a;
			11'h00e: dataout<=36'h7d1806c6f;
			11'h00f: dataout<=36'ha79368dd1;
			11'h010: dataout<=36'h484825974;
			11'h011: dataout<=36'h88b18b973;
			11'h012: dataout<=36'h7ca487471;
			11'h013: dataout<=36'ha99268658;
			11'h014: dataout<=36'h48d825b01;
			11'h015: dataout<=36'h8834cb458;
			11'h016: dataout<=36'h7c28c7c68;
			11'h017: dataout<=36'hab9ba7f0c;
			11'h018: dataout<=36'h4967e5c91;
			11'h019: dataout<=36'h87bb0af37;
			11'h01a: dataout<=36'h7ba54845a;
			11'h01b: dataout<=36'hadaea77ed;
			11'h01c: dataout<=36'h49f6e5e23;
			11'h01d: dataout<=36'h87450aa13;
			11'h01e: dataout<=36'h7b1a08c40;
			11'h01f: dataout<=36'hafcb670fc;
			11'h020: dataout<=36'h4a8565fb9;
			11'h021: dataout<=36'h86d28a4e8;
			11'h022: dataout<=36'h7a864941f;
			11'h023: dataout<=36'hb1f166a3a;
			11'h024: dataout<=36'h4b1366152;
			11'h025: dataout<=36'h866389fb8;
			11'h026: dataout<=36'h79ea49bf4;
			11'h027: dataout<=36'hb420a63a6;
			11'h028: dataout<=36'h4ba0e62ee;
			11'h029: dataout<=36'h85f809a84;
			11'h02a: dataout<=36'h79468a3bf;
			11'h02b: dataout<=36'hb658a5d43;
			11'h02c: dataout<=36'h4c2da648d;
			11'h02d: dataout<=36'h85908954c;
			11'h02e: dataout<=36'h789a8ab7d;
			11'h02f: dataout<=36'hb89925711;
			11'h030: dataout<=36'h4cba2662f;
			11'h031: dataout<=36'h852bc900e;
			11'h032: dataout<=36'h77e70b335;
			11'h033: dataout<=36'hbae225110;
			11'h034: dataout<=36'h4d45e67d4;
			11'h035: dataout<=36'h84cb48acd;
			11'h036: dataout<=36'h772b4badd;
			11'h037: dataout<=36'hbd3324b42;
			11'h038: dataout<=36'h4dd0e697c;
			11'h039: dataout<=36'h846e88588;
			11'h03a: dataout<=36'h76678c277;
			11'h03b: dataout<=36'hbf8be45a7;
			11'h03c: dataout<=36'h4e5ba6b27;
			11'h03d: dataout<=36'h8414c803f;
			11'h03e: dataout<=36'h759c8ca08;
			11'h03f: dataout<=36'hc1ec2403f;
			11'h040: dataout<=36'h4ee5a6cd5;
			11'h041: dataout<=36'h83bf47af2;
			11'h042: dataout<=36'h74c94d18a;
			11'h043: dataout<=36'hc453e3b0c;
			11'h044: dataout<=36'h4f6f26e86;
			11'h045: dataout<=36'h836d075a1;
			11'h046: dataout<=36'h73ee8d8ff;
			11'h047: dataout<=36'hc6c26360d;
			11'h048: dataout<=36'h4ff82703a;
			11'h049: dataout<=36'h831e4704c;
			11'h04a: dataout<=36'h730c4e067;
			11'h04b: dataout<=36'hc937a3144;
			11'h04c: dataout<=36'h5080671f0;
			11'h04d: dataout<=36'h82d346af6;
			11'h04e: dataout<=36'h7222ce7bd;
			11'h04f: dataout<=36'hcbb362cb1;
			11'h050: dataout<=36'h5108273aa;
			11'h051: dataout<=36'h828c0659b;
			11'h052: dataout<=36'h71314ef07;
			11'h053: dataout<=36'hce3522855;
			11'h054: dataout<=36'h518f27566;
			11'h055: dataout<=36'h824886040;
			11'h056: dataout<=36'h70390f63d;
			11'h057: dataout<=36'hd0bca2430;
			11'h058: dataout<=36'h5215a7726;
			11'h059: dataout<=36'h8208c5adf;
			11'h05a: dataout<=36'h6f388fd65;
			11'h05b: dataout<=36'hd349a2042;
			11'h05c: dataout<=36'h529ba78e8;
			11'h05d: dataout<=36'h81cc8557c;
			11'h05e: dataout<=36'h6e311047e;
			11'h05f: dataout<=36'hd5dbe1c8c;
			11'h060: dataout<=36'h532127aad;
			11'h061: dataout<=36'h819385016;
			11'h062: dataout<=36'h6d2290b87;
			11'h063: dataout<=36'hd8732190f;
			11'h064: dataout<=36'h53a5a7c75;
			11'h065: dataout<=36'h815f04ab0;
			11'h066: dataout<=36'h6c0cd1279;
			11'h067: dataout<=36'hdb0ee15ca;
			11'h068: dataout<=36'h5429e7e40;
			11'h069: dataout<=36'h812dc4545;
			11'h06a: dataout<=36'h6aef9195d;
			11'h06b: dataout<=36'hddaf212bf;
			11'h06c: dataout<=36'h54ad6800d;
			11'h06d: dataout<=36'h810003fda;
			11'h06e: dataout<=36'h69cc1202e;
			11'h06f: dataout<=36'he05360fed;
			11'h070: dataout<=36'h5530681de;
			11'h071: dataout<=36'h80d683a6b;
			11'h072: dataout<=36'h68a0926ed;
			11'h073: dataout<=36'he2fb20d56;
			11'h074: dataout<=36'h55b2a83b1;
			11'h075: dataout<=36'h80b0434fc;
			11'h076: dataout<=36'h676f12d97;
			11'h077: dataout<=36'he5a660af8;
			11'h078: dataout<=36'h563428587;
			11'h079: dataout<=36'h808e42f8c;
			11'h07a: dataout<=36'h66365342c;
			11'h07b: dataout<=36'he854a08d5;
			11'h07c: dataout<=36'h56b52875f;
			11'h07d: dataout<=36'h806f42a1b;
			11'h07e: dataout<=36'h64f7d3aae;
			11'h07f: dataout<=36'heb05e06ed;
			11'h080: dataout<=36'h5735a893b;
			11'h081: dataout<=36'h8054824a6;
			11'h082: dataout<=36'h63b15411d;
			11'h083: dataout<=36'hedb960540;
			11'h084: dataout<=36'h57b568b19;
			11'h085: dataout<=36'h803d41f31;
			11'h086: dataout<=36'h626514776;
			11'h087: dataout<=36'hf06ee03cd;
			11'h088: dataout<=36'h583468cfa;
			11'h089: dataout<=36'h802a019bc;
			11'h08a: dataout<=36'h611214db8;
			11'h08b: dataout<=36'hf32660297;
			11'h08c: dataout<=36'h58b2e8ede;
			11'h08d: dataout<=36'h801a41445;
			11'h08e: dataout<=36'h5fb8953e6;
			11'h08f: dataout<=36'hf5df6019b;
			11'h090: dataout<=36'h5930a90c4;
			11'h091: dataout<=36'h800e40ecf;
			11'h092: dataout<=36'h5e59159fc;
			11'h093: dataout<=36'hf899a00dc;
			11'h094: dataout<=36'h59ade92ad;
			11'h095: dataout<=36'h800600958;
			11'h096: dataout<=36'h5cf355ffc;
			11'h097: dataout<=36'hfb54a0058;
			11'h098: dataout<=36'h5a2a69498;
			11'h099: dataout<=36'h8001403e1;
			11'h09a: dataout<=36'h5b87d65e5;
			11'h09b: dataout<=36'hfe1020010;
			11'h09c: dataout<=36'h5aa629687;
			11'h09d: dataout<=36'h8000ffe69;
			11'h09e: dataout<=36'h5a1596bb6;
			11'h09f: dataout<=36'h00cbe0003;
			11'h0a0: dataout<=36'h5b2169878;
			11'h0a1: dataout<=36'h8003ff8f1;
			11'h0a2: dataout<=36'h589d97170;
			11'h0a3: dataout<=36'h038760032;
			11'h0a4: dataout<=36'h5b9be9a6b;
			11'h0a5: dataout<=36'h800a7f37a;
			11'h0a6: dataout<=36'h572057711;
			11'h0a7: dataout<=36'h0642e009d;
			11'h0a8: dataout<=36'h5c15e9c61;
			11'h0a9: dataout<=36'h80147ee03;
			11'h0aa: dataout<=36'h559d57c9c;
			11'h0ab: dataout<=36'h08fd60144;
			11'h0ac: dataout<=36'h5c8ee9e5a;
			11'h0ad: dataout<=36'h8022fe88d;
			11'h0ae: dataout<=36'h541458209;
			11'h0af: dataout<=36'h0bb6e0227;
			11'h0b0: dataout<=36'h5d076a056;
			11'h0b1: dataout<=36'h80353e316;
			11'h0b2: dataout<=36'h52851875f;
			11'h0b3: dataout<=36'h0e6ee0344;
			11'h0b4: dataout<=36'h5d7f6a253;
			11'h0b5: dataout<=36'h804a3dda2;
			11'h0b6: dataout<=36'h50f218c9e;
			11'h0b7: dataout<=36'h11256049e;
			11'h0b8: dataout<=36'h5df66a454;
			11'h0b9: dataout<=36'h8063fd82e;
			11'h0ba: dataout<=36'h4f58591bf;
			11'h0bb: dataout<=36'h13d9e0632;
			11'h0bc: dataout<=36'h5e6cea657;
			11'h0bd: dataout<=36'h8080fd2bb;
			11'h0be: dataout<=36'h4dba196c8;
			11'h0bf: dataout<=36'h168c20802;
			11'h0c0: dataout<=36'h5ee2aa85c;
			11'h0c1: dataout<=36'h80a1bcd4a;
			11'h0c2: dataout<=36'h4c1699bb5;
			11'h0c3: dataout<=36'h193ba0a0c;
			11'h0c4: dataout<=36'h5f57eaa64;
			11'h0c5: dataout<=36'h80c5fc7d9;
			11'h0c6: dataout<=36'h4a6e1a089;
			11'h0c7: dataout<=36'h1be820c52;
			11'h0c8: dataout<=36'h5fcc2ac6f;
			11'h0c9: dataout<=36'h80ee7c26b;
			11'h0ca: dataout<=36'h48c09a53f;
			11'h0cb: dataout<=36'h1e9160ed1;
			11'h0cc: dataout<=36'h603feae7c;
			11'h0cd: dataout<=36'h811a7bcfe;
			11'h0ce: dataout<=36'h470e1a9db;
			11'h0cf: dataout<=36'h21372118a;
			11'h0d0: dataout<=36'h60b2eb08b;
			11'h0d1: dataout<=36'h8149bb794;
			11'h0d2: dataout<=36'h4557dae5b;
			11'h0d3: dataout<=36'h23d92147e;
			11'h0d4: dataout<=36'h61252b29d;
			11'h0d5: dataout<=36'h817d3b22c;
			11'h0d6: dataout<=36'h439c5b2bd;
			11'h0d7: dataout<=36'h2676a17aa;
			11'h0d8: dataout<=36'h6196ab4b2;
			11'h0d9: dataout<=36'h81b4bacc5;
			11'h0da: dataout<=36'h41dbdb703;
			11'h0db: dataout<=36'h290fe1b10;
			11'h0dc: dataout<=36'h6207ab6c8;
			11'h0dd: dataout<=36'h81eefa761;
			11'h0de: dataout<=36'h40181bb2f;
			11'h0df: dataout<=36'h2ba461eae;
			11'h0e0: dataout<=36'h6277ab8e2;
			11'h0e1: dataout<=36'h822dba200;
			11'h0e2: dataout<=36'h3e4f5bf3a;
			11'h0e3: dataout<=36'h2e33a2285;
			11'h0e4: dataout<=36'h62e72bafd;
			11'h0e5: dataout<=36'h826f79ca2;
			11'h0e6: dataout<=36'h3c831c32a;
			11'h0e7: dataout<=36'h30bd62693;
			11'h0e8: dataout<=36'h6355ebd1b;
			11'h0e9: dataout<=36'h82b539746;
			11'h0ea: dataout<=36'h3ab29c6fc;
			11'h0eb: dataout<=36'h3341a2ad8;
			11'h0ec: dataout<=36'h63c3abf3b;
			11'h0ed: dataout<=36'h82feb91ef;
			11'h0ee: dataout<=36'h38de9caae;
			11'h0ef: dataout<=36'h35bfe2f55;
			11'h0f0: dataout<=36'h6430ec15e;
			11'h0f1: dataout<=36'h834bf8c99;
			11'h0f2: dataout<=36'h37061ce43;
			11'h0f3: dataout<=36'h3837e3407;
			11'h0f4: dataout<=36'h649d6c383;
			11'h0f5: dataout<=36'h839cb8747;
			11'h0f6: dataout<=36'h352a9d1ba;
			11'h0f7: dataout<=36'h3aa9238ef;
			11'h0f8: dataout<=36'h65096c5aa;
			11'h0f9: dataout<=36'h83f0b81f8;
			11'h0fa: dataout<=36'h334b5d515;
			11'h0fb: dataout<=36'h3d13e3e0d;
			11'h0fc: dataout<=36'h65746c7d4;
			11'h0fd: dataout<=36'h8448b7cad;
			11'h0fe: dataout<=36'h31689d84f;
			11'h0ff: dataout<=36'h3f772435f;
			11'h100: dataout<=36'h65deaca00;
			11'h101: dataout<=36'h84a477766;
			11'h102: dataout<=36'h2f829db69;
			11'h103: dataout<=36'h41d3248e4;
			11'h104: dataout<=36'h66482cc2e;
			11'h105: dataout<=36'h8503b7224;
			11'h106: dataout<=36'h2d99dde64;
			11'h107: dataout<=36'h442764e9d;
			11'h108: dataout<=36'h66b0ece5e;
			11'h109: dataout<=36'h856676ce6;
			11'h10a: dataout<=36'h2bae5e13f;
			11'h10b: dataout<=36'h4673e5489;
			11'h10c: dataout<=36'h67192d091;
			11'h10d: dataout<=36'h85ccb67aa;
			11'h10e: dataout<=36'h29bf1e3fe;
			11'h10f: dataout<=36'h48b7e5aa7;
			11'h110: dataout<=36'h67806d2c5;
			11'h111: dataout<=36'h863636275;
			11'h112: dataout<=36'h27ce5e69b;
			11'h113: dataout<=36'h4af3a60f5;
			11'h114: dataout<=36'h67e6ed4fc;
			11'h115: dataout<=36'h86a3b5d44;
			11'h116: dataout<=36'h25da1e917;
			11'h117: dataout<=36'h4d2666775;
			11'h118: dataout<=36'h684cad736;
			11'h119: dataout<=36'h871535817;
			11'h11a: dataout<=36'h23e31eb72;
			11'h11b: dataout<=36'h4f5066e24;
			11'h11c: dataout<=36'h68b1ed971;
			11'h11d: dataout<=36'h8789352ee;
			11'h11e: dataout<=36'h21ea1edb2;
			11'h11f: dataout<=36'h5170e7502;
			11'h120: dataout<=36'h69162dbae;
			11'h121: dataout<=36'h880134dcc;
			11'h122: dataout<=36'h1fef1efce;
			11'h123: dataout<=36'h538827c0e;
			11'h124: dataout<=36'h6979addee;
			11'h125: dataout<=36'h887cf48ae;
			11'h126: dataout<=36'h1df19f1c9;
			11'h127: dataout<=36'h559568347;
			11'h128: dataout<=36'h69dc6e030;
			11'h129: dataout<=36'h88fbf4395;
			11'h12a: dataout<=36'h1bf21f3a4;
			11'h12b: dataout<=36'h5798a8aad;
			11'h12c: dataout<=36'h6a3e2e274;
			11'h12d: dataout<=36'h897eb3e84;
			11'h12e: dataout<=36'h19f15f55b;
			11'h12f: dataout<=36'h5991e923e;
			11'h130: dataout<=36'h6a9f6e4b9;
			11'h131: dataout<=36'h8a0433978;
			11'h132: dataout<=36'h17ef1f6f6;
			11'h133: dataout<=36'h5b80a99fa;
			11'h134: dataout<=36'h6affee701;
			11'h135: dataout<=36'h8a8db3470;
			11'h136: dataout<=36'h15ea9f86e;
			11'h137: dataout<=36'h5d646a1e0;
			11'h138: dataout<=36'h6b5f6e94b;
			11'h139: dataout<=36'h8b1ab2f6f;
			11'h13a: dataout<=36'h13e49f9c4;
			11'h13b: dataout<=36'h5f3daa9ef;
			11'h13c: dataout<=36'h6bbe6eb98;
			11'h13d: dataout<=36'h8baaf2a72;
			11'h13e: dataout<=36'h11dcdfafb;
			11'h13f: dataout<=36'h610bab225;
			11'h140: dataout<=36'h6c1c6ede6;
			11'h141: dataout<=36'h8c3eb257e;
			11'h142: dataout<=36'h0fd4dfc0e;
			11'h143: dataout<=36'h62ce2ba83;
			11'h144: dataout<=36'h6c79af036;
			11'h145: dataout<=36'h8cd5b208f;
			11'h146: dataout<=36'h0dcb5fd02;
			11'h147: dataout<=36'h64852c307;
			11'h148: dataout<=36'h6cd62f288;
			11'h149: dataout<=36'h8d6ff1ba7;
			11'h14a: dataout<=36'h0bc15fdd4;
			11'h14b: dataout<=36'h6630acbaf;
			11'h14c: dataout<=36'h6d31ef4dc;
			11'h14d: dataout<=36'h8e0db16c5;
			11'h14e: dataout<=36'h09b61fe84;
			11'h14f: dataout<=36'h67d02d47c;
			11'h150: dataout<=36'h6d8caf732;
			11'h151: dataout<=36'h8eaef11ec;
			11'h152: dataout<=36'h07aadff11;
			11'h153: dataout<=36'h69636dd6b;
			11'h154: dataout<=36'h6de6ef98a;
			11'h155: dataout<=36'h8f5330d17;
			11'h156: dataout<=36'h059e5ff7f;
			11'h157: dataout<=36'h6aea6e67d;
			11'h158: dataout<=36'h6e402fbe4;
			11'h159: dataout<=36'h8ffaf084b;
			11'h15a: dataout<=36'h0391dffca;
			11'h15b: dataout<=36'h6c64eefaf;
			11'h15c: dataout<=36'h6e98afe3f;
			11'h15d: dataout<=36'h90a570386;
			11'h15e: dataout<=36'h01855fff5;
			11'h15f: dataout<=36'h6dd2af902;
			11'h160: dataout<=36'h6ef03009d;
			11'h161: dataout<=36'h9153efec9;
			11'h162: dataout<=36'hff789fffb;
			11'h163: dataout<=36'h6f33b0273;
			11'h164: dataout<=36'h6f47302fc;
			11'h165: dataout<=36'h9204efa12;
			11'h166: dataout<=36'hfd6bdffe4;
			11'h167: dataout<=36'h7087f0c01;
			11'h168: dataout<=36'h6f9d3055e;
			11'h169: dataout<=36'h92b9ef563;
			11'h16a: dataout<=36'hfb5edffa7;
			11'h16b: dataout<=36'h71ceb15ac;
			11'h16c: dataout<=36'h6ff2707c1;
			11'h16d: dataout<=36'h9371af0bc;
			11'h16e: dataout<=36'hf9529ff4b;
			11'h16f: dataout<=36'h730871f73;
			11'h170: dataout<=36'h7046f0a26;
			11'h171: dataout<=36'h942caec1c;
			11'h172: dataout<=36'hf7465fecd;
			11'h173: dataout<=36'h743472953;
			11'h174: dataout<=36'h709a70c8d;
			11'h175: dataout<=36'h94eaee786;
			11'h176: dataout<=36'hf53b5fe2c;
			11'h177: dataout<=36'h75533334d;
			11'h178: dataout<=36'h70ed30ef5;
			11'h179: dataout<=36'h95abee2f8;
			11'h17a: dataout<=36'hf3311fd6b;
			11'h17b: dataout<=36'h766433d5e;
			11'h17c: dataout<=36'h713f3115f;
			11'h17d: dataout<=36'h96702de71;
			11'h17e: dataout<=36'hf1275fc89;
			11'h17f: dataout<=36'h776734787;
			11'h180: dataout<=36'h7190313cb;
			11'h181: dataout<=36'h9737ad9f4;
			11'h182: dataout<=36'hef1edfb84;
			11'h183: dataout<=36'h785c751c5;
			11'h184: dataout<=36'h71e0b1639;
			11'h185: dataout<=36'h98022d57d;
			11'h186: dataout<=36'hed169fa5f;
			11'h187: dataout<=36'h794375c17;
			11'h188: dataout<=36'h7230318a9;
			11'h189: dataout<=36'h98cfed10f;
			11'h18a: dataout<=36'heb0f9f918;
			11'h18b: dataout<=36'h7a1c7667c;
			11'h18c: dataout<=36'h727eb1b1a;
			11'h18d: dataout<=36'h99a06ccad;
			11'h18e: dataout<=36'he90b1f7af;
			11'h18f: dataout<=36'h7ae7370f3;
			11'h190: dataout<=36'h72cc71d8d;
			11'h191: dataout<=36'h9a742c852;
			11'h192: dataout<=36'he7075f625;
			11'h193: dataout<=36'h7ba377b7b;
			11'h194: dataout<=36'h731972001;
			11'h195: dataout<=36'h9b4a2c400;
			11'h196: dataout<=36'he5059f47d;
			11'h197: dataout<=36'h7c5178613;
			11'h198: dataout<=36'h7365b2277;
			11'h199: dataout<=36'h9c23abfb7;
			11'h19a: dataout<=36'he3055f2b3;
			11'h19b: dataout<=36'h7cf0b90b8;
			11'h19c: dataout<=36'h73b0f24ef;
			11'h19d: dataout<=36'h9d002bb77;
			11'h19e: dataout<=36'he106df0c6;
			11'h19f: dataout<=36'h7d8179b6b;
			11'h1a0: dataout<=36'h73fb32768;
			11'h1a1: dataout<=36'h9ddf2b743;
			11'h1a2: dataout<=36'hdf0b5eeba;
			11'h1a3: dataout<=36'h7e03ba62a;
			11'h1a4: dataout<=36'h7444f29e3;
			11'h1a5: dataout<=36'h9ec16b316;
			11'h1a6: dataout<=36'hdd10dec8d;
			11'h1a7: dataout<=36'h7e773b0f2;
			11'h1a8: dataout<=36'h748db2c60;
			11'h1a9: dataout<=36'h9fa66aef3;
			11'h1aa: dataout<=36'hdb18dea40;
			11'h1ab: dataout<=36'h7edbbbbc5;
			11'h1ac: dataout<=36'h74d572ede;
			11'h1ad: dataout<=36'ha08e6aadb;
			11'h1ae: dataout<=36'hd9239e7d1;
			11'h1af: dataout<=36'h7f31bc69f;
			11'h1b0: dataout<=36'h751c7315d;
			11'h1b1: dataout<=36'ha178aa6cd;
			11'h1b2: dataout<=36'hd7311e545;
			11'h1b3: dataout<=36'h7f78bd17f;
			11'h1b4: dataout<=36'h7562b33de;
			11'h1b5: dataout<=36'ha265ea2c8;
			11'h1b6: dataout<=36'hd5411e298;
			11'h1b7: dataout<=36'h7fb0bdc66;
			11'h1b8: dataout<=36'h75a833661;
			11'h1b9: dataout<=36'ha355e9ecc;
			11'h1ba: dataout<=36'hd3531dfcc;
			11'h1bb: dataout<=36'h7fd9fe750;
			11'h1bc: dataout<=36'h75ec738e5;
			11'h1bd: dataout<=36'ha448e9ade;
			11'h1be: dataout<=36'hd1695dcdd;
			11'h1bf: dataout<=36'h7ff43f23d;
			11'h1c0: dataout<=36'h763033b6a;
			11'h1c1: dataout<=36'ha53de96f7;
			11'h1c2: dataout<=36'hcf81dd9d4;
			11'h1c3: dataout<=36'h7fff7fd2c;
			11'h1c4: dataout<=36'h7672f3df1;
			11'h1c5: dataout<=36'ha6362931c;
			11'h1c6: dataout<=36'hcd9d9d6a8;
			11'h1c7: dataout<=36'h7ffbc081a;
			11'h1c8: dataout<=36'h76b4b4079;
			11'h1c9: dataout<=36'ha730a8f4d;
			11'h1ca: dataout<=36'hcbbd5d35e;
			11'h1cb: dataout<=36'h7fe941309;
			11'h1cc: dataout<=36'h76f5b4303;
			11'h1cd: dataout<=36'ha82e28b87;
			11'h1ce: dataout<=36'hc9dfdcff5;
			11'h1cf: dataout<=36'h7fc7c1df5;
			11'h1d0: dataout<=36'h7735f458e;
			11'h1d1: dataout<=36'ha92de87cb;
			11'h1d2: dataout<=36'hc8059cc6f;
			11'h1d3: dataout<=36'h7f97428dd;
			11'h1d4: dataout<=36'h77753481b;
			11'h1d5: dataout<=36'haa306841b;
			11'h1d6: dataout<=36'hc62f5c8c9;
			11'h1d7: dataout<=36'h7f58033c1;
			11'h1d8: dataout<=36'h77b3b4aa8;
			11'h1d9: dataout<=36'hab34e8076;
			11'h1da: dataout<=36'hc45d1c508;
			11'h1db: dataout<=36'h7f09c3e9f;
			11'h1dc: dataout<=36'h77f134d38;
			11'h1dd: dataout<=36'hac3ca7cdc;
			11'h1de: dataout<=36'hc28e5c125;
			11'h1df: dataout<=36'h7eacc4975;
			11'h1e0: dataout<=36'h782db4fc8;
			11'h1e1: dataout<=36'had4667950;
			11'h1e2: dataout<=36'hc0c49bd26;
			11'h1e3: dataout<=36'h7e4105443;
			11'h1e4: dataout<=36'h7869b525a;
			11'h1e5: dataout<=36'hae52a75cb;
			11'h1e6: dataout<=36'hbefddb90b;
			11'h1e7: dataout<=36'h7dc685f07;
			11'h1e8: dataout<=36'h78a4754ed;
			11'h1e9: dataout<=36'haf6127255;
			11'h1ea: dataout<=36'hbd3c5b4d2;
			11'h1eb: dataout<=36'h7d3d469c0;
			11'h1ec: dataout<=36'h78de75781;
			11'h1ed: dataout<=36'hb07226ee9;
			11'h1ee: dataout<=36'hbb7e9b07c;
			11'h1ef: dataout<=36'h7ca58746c;
			11'h1f0: dataout<=36'h7917b5a16;
			11'h1f1: dataout<=36'hb18526b89;
			11'h1f2: dataout<=36'hb9c59ac0c;
			11'h1f3: dataout<=36'h7bff07f0b;
			11'h1f4: dataout<=36'h794ff5cad;
			11'h1f5: dataout<=36'hb29ae6834;
			11'h1f6: dataout<=36'hb810da77d;
			11'h1f7: dataout<=36'h7b4a4899b;
			11'h1f8: dataout<=36'h798735f45;
			11'h1f9: dataout<=36'hb3b2e64ed;
			11'h1fa: dataout<=36'hb6615a2d2;
			11'h1fb: dataout<=36'h7a870941b;
			11'h1fc: dataout<=36'h79bdb61de;
			11'h1fd: dataout<=36'hb4cce61b0;
			11'h1fe: dataout<=36'hb4b659e0d;
			11'h1ff: dataout<=36'h79b549e8a;
			11'h200: dataout<=36'h79f376478;
			11'h201: dataout<=36'hb5e8e5e7f;
			11'h202: dataout<=36'hb3101992f;
			11'h203: dataout<=36'h78d58a8e6;
			11'h204: dataout<=36'h7a27f6713;
			11'h205: dataout<=36'hb70725b5c;
			11'h206: dataout<=36'hb16fd9433;
			11'h207: dataout<=36'h77e7cb32f;
			11'h208: dataout<=36'h7a5bf69b0;
			11'h209: dataout<=36'hb827e5843;
			11'h20a: dataout<=36'hafd358f1d;
			11'h20b: dataout<=36'h76ebcbd63;
			11'h20c: dataout<=36'h7a8eb6c4d;
			11'h20d: dataout<=36'hb94a65539;
			11'h20e: dataout<=36'hae3d589ed;
			11'h20f: dataout<=36'h75e20c780;
			11'h210: dataout<=36'h7ac0b6eec;
			11'h211: dataout<=36'hba6f6523a;
			11'h212: dataout<=36'hacac184a2;
			11'h213: dataout<=36'h74ca8d186;
			11'h214: dataout<=36'h7af1f718c;
			11'h215: dataout<=36'hbb9624f47;
			11'h216: dataout<=36'hab2057f3e;
			11'h217: dataout<=36'h73a54db74;
			11'h218: dataout<=36'h7b223742c;
			11'h219: dataout<=36'hbcbea4c61;
			11'h21a: dataout<=36'ha99a579c3;
			11'h21b: dataout<=36'h72728e548;
			11'h21c: dataout<=36'h7b51776ce;
			11'h21d: dataout<=36'hbde964988;
			11'h21e: dataout<=36'ha819d742d;
			11'h21f: dataout<=36'h71328ef01;
			11'h220: dataout<=36'h7b7ff7971;
			11'h221: dataout<=36'hbf16246bb;
			11'h222: dataout<=36'ha69ed6e7f;
			11'h223: dataout<=36'h6fe54f89f;
			11'h224: dataout<=36'h7bad77c14;
			11'h225: dataout<=36'hc044643fd;
			11'h226: dataout<=36'ha52a968ba;
			11'h227: dataout<=36'h6e8b1021f;
			11'h228: dataout<=36'h7bd9f7eb9;
			11'h229: dataout<=36'hc174e414b;
			11'h22a: dataout<=36'ha3bc162db;
			11'h22b: dataout<=36'h6d23d0b81;
			11'h22c: dataout<=36'h7c05b815f;
			11'h22d: dataout<=36'hc2a723ea5;
			11'h22e: dataout<=36'ha25315ce6;
			11'h22f: dataout<=36'h6bafd14c4;
			11'h230: dataout<=36'h7c30b8405;
			11'h231: dataout<=36'hc3dae3c0c;
			11'h232: dataout<=36'ha0f0556dc;
			11'h233: dataout<=36'h6a2f11de7;
			11'h234: dataout<=36'h7c5a786ad;
			11'h235: dataout<=36'hc510e3982;
			11'h236: dataout<=36'h9f94150b8;
			11'h237: dataout<=36'h68a2526e9;
			11'h238: dataout<=36'h7c8378955;
			11'h239: dataout<=36'hc64863704;
			11'h23a: dataout<=36'h9e3e14a7f;
			11'h23b: dataout<=36'h670912fc7;
			11'h23c: dataout<=36'h7cabb8bfe;
			11'h23d: dataout<=36'hc78163493;
			11'h23e: dataout<=36'h9cee54432;
			11'h23f: dataout<=36'h6563d3883;
			11'h240: dataout<=36'h7cd2b8ea8;
			11'h241: dataout<=36'hc8bc23231;
			11'h242: dataout<=36'h9ba5d3dcf;
			11'h243: dataout<=36'h63b2d411a;
			11'h244: dataout<=36'h7cf8f9153;
			11'h245: dataout<=36'hc9f8a2fdc;
			11'h246: dataout<=36'h9a6353756;
			11'h247: dataout<=36'h61f61498b;
			11'h248: dataout<=36'h7d1e793ff;
			11'h249: dataout<=36'hcb36a2d93;
			11'h24a: dataout<=36'h9927130c9;
			11'h24b: dataout<=36'h602e151d6;
			11'h24c: dataout<=36'h7d42f96ab;
			11'h24d: dataout<=36'hcc75e2b58;
			11'h24e: dataout<=36'h97f212a2a;
			11'h24f: dataout<=36'h5e5a959fa;
			11'h250: dataout<=36'h7d6679958;
			11'h251: dataout<=36'hcdb6e292c;
			11'h252: dataout<=36'h96c412375;
			11'h253: dataout<=36'h5c7c561f5;
			11'h254: dataout<=36'h7d88f9c06;
			11'h255: dataout<=36'hcef96270e;
			11'h256: dataout<=36'h959d11cad;
			11'h257: dataout<=36'h5a93169c7;
			11'h258: dataout<=36'h7daab9eb5;
			11'h259: dataout<=36'hd03da24fc;
			11'h25a: dataout<=36'h947c515d2;
			11'h25b: dataout<=36'h589f5716e;
			11'h25c: dataout<=36'h7dcb7a165;
			11'h25d: dataout<=36'hd183222f9;
			11'h25e: dataout<=36'h936310ee4;
			11'h25f: dataout<=36'h56a1578eb;
			11'h260: dataout<=36'h7deb7a415;
			11'h261: dataout<=36'hd2c9a2102;
			11'h262: dataout<=36'h9250907e7;
			11'h263: dataout<=36'h54991803b;
			11'h264: dataout<=36'h7e0a7a6c6;
			11'h265: dataout<=36'hd411e1f1a;
			11'h266: dataout<=36'h9145500d6;
			11'h267: dataout<=36'h52871875f;
			11'h268: dataout<=36'h7e287a977;
			11'h269: dataout<=36'hd55ae1d42;
			11'h26a: dataout<=36'h90420f9b7;
			11'h26b: dataout<=36'h506b58e54;
			11'h26c: dataout<=36'h7e457ac29;
			11'h26d: dataout<=36'hd6a561b77;
			11'h26e: dataout<=36'h8f460f286;
			11'h26f: dataout<=36'h4e461951c;
			11'h270: dataout<=36'h7e61baedc;
			11'h271: dataout<=36'hd7f1619b9;
			11'h272: dataout<=36'h8e50ceb44;
			11'h273: dataout<=36'h4c17d9bb4;
			11'h274: dataout<=36'h7e7cfb18f;
			11'h275: dataout<=36'hd93e2180b;
			11'h276: dataout<=36'h8d638e3f5;
			11'h277: dataout<=36'h49e0da21c;
			11'h278: dataout<=36'h7e973b443;
			11'h279: dataout<=36'hda8c6166b;
			11'h27a: dataout<=36'h8c7dcdc94;
			11'h27b: dataout<=36'h47a11a853;
			11'h27c: dataout<=36'h7eb0bb6f7;
			11'h27d: dataout<=36'hdbdb214d8;
			11'h27e: dataout<=36'h8b9f8d529;
			11'h27f: dataout<=36'h4558dae58;
			11'h280: dataout<=36'h7ec93b9ac;
			11'h281: dataout<=36'hdd2b61354;
			11'h282: dataout<=36'h8ac8ccdad;
			11'h283: dataout<=36'h43089b42c;
			11'h284: dataout<=36'h7ee0bbc62;
			11'h285: dataout<=36'hde7ce11de;
			11'h286: dataout<=36'h89f98c622;
			11'h287: dataout<=36'h40b09b9cc;
			11'h288: dataout<=36'h7ef77bf17;
			11'h289: dataout<=36'hdfcea1077;
			11'h28a: dataout<=36'h89328be8e;
			11'h28b: dataout<=36'h3e511bf39;
			11'h28c: dataout<=36'h7f0d3c1ce;
			11'h28d: dataout<=36'he12220f1d;
			11'h28e: dataout<=36'h88728b6e9;
			11'h28f: dataout<=36'h3bea1c472;
			11'h290: dataout<=36'h7f21fc485;
			11'h291: dataout<=36'he27620dd3;
			11'h292: dataout<=36'h87bb4af3a;
			11'h293: dataout<=36'h397c5c975;
			11'h294: dataout<=36'h7f35bc73c;
			11'h295: dataout<=36'he3cae0c99;
			11'h296: dataout<=36'h870c0a781;
			11'h297: dataout<=36'h37079ce44;
			11'h298: dataout<=36'h7f48bc9f4;
			11'h299: dataout<=36'he520a0b6b;
			11'h29a: dataout<=36'h866409fbb;
			11'h29b: dataout<=36'h348c9d2dc;
			11'h29c: dataout<=36'h7f5abccac;
			11'h29d: dataout<=36'he67720a4c;
			11'h29e: dataout<=36'h85c4497eb;
			11'h29f: dataout<=36'h320b9d73e;
			11'h2a0: dataout<=36'h7f6bbcf64;
			11'h2a1: dataout<=36'he7ce2093d;
			11'h2a2: dataout<=36'h852cc9013;
			11'h2a3: dataout<=36'h2f849db69;
			11'h2a4: dataout<=36'h7f7bfd21d;
			11'h2a5: dataout<=36'he9262083b;
			11'h2a6: dataout<=36'h849cc882f;
			11'h2a7: dataout<=36'h2cf81df5c;
			11'h2a8: dataout<=36'h7f8b3d4d6;
			11'h2a9: dataout<=36'hea7ea0748;
			11'h2aa: dataout<=36'h841508044;
			11'h2ab: dataout<=36'h2a665e318;
			11'h2ac: dataout<=36'h7f997d790;
			11'h2ad: dataout<=36'hebd820665;
			11'h2ae: dataout<=36'h83960784e;
			11'h2af: dataout<=36'h27cf9e69b;
			11'h2b0: dataout<=36'h7fa6bda4a;
			11'h2b1: dataout<=36'hed3220591;
			11'h2b2: dataout<=36'h831f07050;
			11'h2b3: dataout<=36'h25341e9e5;
			11'h2b4: dataout<=36'h7fb33dd04;
			11'h2b5: dataout<=36'hee8ca04ca;
			11'h2b6: dataout<=36'h82afc684c;
			11'h2b7: dataout<=36'h22945ecf6;
			11'h2b8: dataout<=36'h7fbebdfbe;
			11'h2b9: dataout<=36'hefe720412;
			11'h2ba: dataout<=36'h8248c6043;
			11'h2bb: dataout<=36'h1ff09efcd;
			11'h2bc: dataout<=36'h7fc93e279;
			11'h2bd: dataout<=36'hf142e036a;
			11'h2be: dataout<=36'h81ea45830;
			11'h2bf: dataout<=36'h1d491f26b;
			11'h2c0: dataout<=36'h7fd2fe533;
			11'h2c1: dataout<=36'hf29e202cf;
			11'h2c2: dataout<=36'h8193c501c;
			11'h2c3: dataout<=36'h1a9e1f4ce;
			11'h2c4: dataout<=36'h7fdbbe7ee;
			11'h2c5: dataout<=36'hf3fa60244;
			11'h2c6: dataout<=36'h8145c4800;
			11'h2c7: dataout<=36'h17f01f6f7;
			11'h2c8: dataout<=36'h7fe37eaa9;
			11'h2c9: dataout<=36'hf556e01c8;
			11'h2ca: dataout<=36'h810003fdf;
			11'h2cb: dataout<=36'h153f5f8e5;
			11'h2cc: dataout<=36'h7fea3ed65;
			11'h2cd: dataout<=36'hf6b42015c;
			11'h2ce: dataout<=36'h80c3037b8;
			11'h2cf: dataout<=36'h128c1fa98;
			11'h2d0: dataout<=36'h7fefff020;
			11'h2d1: dataout<=36'hf810e00fe;
			11'h2d2: dataout<=36'h808e42f91;
			11'h2d3: dataout<=36'h0fd69fc10;
			11'h2d4: dataout<=36'h7ff4ff2dc;
			11'h2d5: dataout<=36'hf96ea00af;
			11'h2d6: dataout<=36'h8061c2763;
			11'h2d7: dataout<=36'h0d1f5fd4d;
			11'h2d8: dataout<=36'h7ff8ff597;
			11'h2d9: dataout<=36'hfacbe006f;
			11'h2da: dataout<=36'h803dc1f36;
			11'h2db: dataout<=36'h0a665fe4e;
			11'h2dc: dataout<=36'h7ffc3f853;
			11'h2dd: dataout<=36'hfc29a003c;
			11'h2de: dataout<=36'h802141705;
			11'h2df: dataout<=36'h07ac5ff14;
			11'h2e0: dataout<=36'h7ffe3fb0f;
			11'h2e1: dataout<=36'hfd87a001b;
			11'h2e2: dataout<=36'h800e80ed2;
			11'h2e3: dataout<=36'h04f15ff9e;
			11'h2e4: dataout<=36'h7fff7fdcb;
			11'h2e5: dataout<=36'hfee5a0007;
			11'h2e6: dataout<=36'h80034069e;
			11'h2e7: dataout<=36'h0235dffec;
			11'h2e8: dataout<=36'h7fff80084;
			11'h2e9: dataout<=36'h004220003;
			11'h2ea: dataout<=36'h80013fe73;
			11'h2eb: dataout<=36'hff7a5fffe;
			11'h2ec: dataout<=36'h7fff00340;
			11'h2ed: dataout<=36'h01a02000c;
			11'h2ee: dataout<=36'h80067f63f;
			11'h2ef: dataout<=36'hfcbe9ffd5;
			11'h2f0: dataout<=36'h7ffd805fc;
			11'h2f1: dataout<=36'h02fe20024;
			11'h2f2: dataout<=36'h80143ee0b;
			11'h2f3: dataout<=36'hfa035ff70;
			11'h2f4: dataout<=36'h7ffac08b8;
			11'h2f5: dataout<=36'h045c2004f;
			11'h2f6: dataout<=36'h802bfe5d9;
			11'h2f7: dataout<=36'hf7489fecf;
			11'h2f8: dataout<=36'h7ff780b73;
			11'h2f9: dataout<=36'h05b960084;
			11'h2fa: dataout<=36'h804a3ddab;
			11'h2fb: dataout<=36'hf48edfdf3;
			11'h2fc: dataout<=36'h7ff300e2f;
			11'h2fd: dataout<=36'h0717200cb;
			11'h2fe: dataout<=36'h8071fd57c;
			11'h2ff: dataout<=36'hf1d69fcdb;
			11'h300: dataout<=36'h7fedc10eb;
			11'h301: dataout<=36'h0874a0120;
			11'h302: dataout<=36'h80a17cd50;
			11'h303: dataout<=36'hef201fb87;
			11'h304: dataout<=36'h7fe7813a6;
			11'h305: dataout<=36'h09d160183;
			11'h306: dataout<=36'h80d97c52a;
			11'h307: dataout<=36'hec6b5f9f9;
			11'h308: dataout<=36'h7fe041661;
			11'h309: dataout<=36'h0b2de01f7;
			11'h30a: dataout<=36'h811a3bd07;
			11'h30b: dataout<=36'he9b8df82f;
			11'h30c: dataout<=36'h7fd84191c;
			11'h30d: dataout<=36'h0c8a60278;
			11'h30e: dataout<=36'h8162fb4e8;
			11'h30f: dataout<=36'he7091f62a;
			11'h310: dataout<=36'h7fcf41bd7;
			11'h311: dataout<=36'h0de660308;
			11'h312: dataout<=36'h81b3bacce;
			11'h313: dataout<=36'he45c5f3eb;
			11'h314: dataout<=36'h7fc541e92;
			11'h315: dataout<=36'h0f42203a7;
			11'h316: dataout<=36'h820d3a4b8;
			11'h317: dataout<=36'he1b29f171;
			11'h318: dataout<=36'h7fba4214c;
			11'h319: dataout<=36'h109d20456;
			11'h31a: dataout<=36'h826f39cab;
			11'h31b: dataout<=36'hdf0c9eebe;
			11'h31c: dataout<=36'h7fae82406;
			11'h31d: dataout<=36'h11f7e0513;
			11'h31e: dataout<=36'h82d8f94a3;
			11'h31f: dataout<=36'hdc6a5ebd0;
			11'h320: dataout<=36'h7fa1826c0;
			11'h321: dataout<=36'h1351e05e0;
			11'h322: dataout<=36'h834bb8ca2;
			11'h323: dataout<=36'hd9cc1e8a9;
			11'h324: dataout<=36'h7f940297a;
			11'h325: dataout<=36'h14abe06b9;
			11'h326: dataout<=36'h83c5784a7;
			11'h327: dataout<=36'hd7329e549;
			11'h328: dataout<=36'h7f8542c33;
			11'h329: dataout<=36'h1604a07a4;
			11'h32a: dataout<=36'h844877cb7;
			11'h32b: dataout<=36'hd49d9e1b1;
			11'h32c: dataout<=36'h7f75c2eec;
			11'h32d: dataout<=36'h175ce089b;
			11'h32e: dataout<=36'h84d2b74ce;
			11'h32f: dataout<=36'hd20dddde0;
			11'h330: dataout<=36'h7f65431a5;
			11'h331: dataout<=36'h18b4e09a2;
			11'h332: dataout<=36'h856576ced;
			11'h333: dataout<=36'hcf835d9d7;
			11'h334: dataout<=36'h7f53c345e;
			11'h335: dataout<=36'h1a0c20ab8;
			11'h336: dataout<=36'h860076515;
			11'h337: dataout<=36'hccfe9d597;
			11'h338: dataout<=36'h7f4183715;
			11'h339: dataout<=36'h1b61e0bdb;
			11'h33a: dataout<=36'h86a2f5d4c;
			11'h33b: dataout<=36'hca7fdd121;
			11'h33c: dataout<=36'h7f2e039cd;
			11'h33d: dataout<=36'h1cb760d10;
			11'h33e: dataout<=36'h874e7558a;
			11'h33f: dataout<=36'hc8071cc73;
			11'h340: dataout<=36'h7f1a03c84;
			11'h341: dataout<=36'h1e0be0e4f;
			11'h342: dataout<=36'h880074dd4;
			11'h343: dataout<=36'hc5951c791;
			11'h344: dataout<=36'h7f04c3f3b;
			11'h345: dataout<=36'h1f5fa0fa0;
			11'h346: dataout<=36'h88bb7462a;
			11'h347: dataout<=36'hc329dc278;
			11'h348: dataout<=36'h7eeec41f1;
			11'h349: dataout<=36'h20b2610fe;
			11'h34a: dataout<=36'h897db3e8c;
			11'h34b: dataout<=36'hc0c5dbd2c;
			11'h34c: dataout<=36'h7ed7c44a7;
			11'h34d: dataout<=36'h22046126b;
			11'h34e: dataout<=36'h8a47f36f9;
			11'h34f: dataout<=36'hbe691b7ab;
			11'h350: dataout<=36'h7ebfc475c;
			11'h351: dataout<=36'h2355213e6;
			11'h352: dataout<=36'h8b19f2f76;
			11'h353: dataout<=36'hbc13db1f7;
			11'h354: dataout<=36'h7ea704a11;
			11'h355: dataout<=36'h24a4e156f;
			11'h356: dataout<=36'h8bf3327ff;
			11'h357: dataout<=36'hb9c6dac10;
			11'h358: dataout<=36'h7e8d44cc5;
			11'h359: dataout<=36'h25f3a1707;
			11'h35a: dataout<=36'h8cd472097;
			11'h35b: dataout<=36'hb781da5f8;
			11'h35c: dataout<=36'h7e7284f79;
			11'h35d: dataout<=36'h2741618ad;
			11'h35e: dataout<=36'h8dbd7193c;
			11'h35f: dataout<=36'hb54559fae;
			11'h360: dataout<=36'h7e56c522c;
			11'h361: dataout<=36'h288de1a63;
			11'h362: dataout<=36'h8eae311f2;
			11'h363: dataout<=36'hb31199934;
			11'h364: dataout<=36'h7e3a454de;
			11'h365: dataout<=36'h29d8e1c25;
			11'h366: dataout<=36'h8fa5b0ab9;
			11'h367: dataout<=36'hb0e6d9289;
			11'h368: dataout<=36'h7e1cc5790;
			11'h369: dataout<=36'h2b22e1df6;
			11'h36a: dataout<=36'h90a4f038e;
			11'h36b: dataout<=36'haec558bb0;
			11'h36c: dataout<=36'h7dfe85a41;
			11'h36d: dataout<=36'h2c6be1fd3;
			11'h36e: dataout<=36'h91aaefc73;
			11'h36f: dataout<=36'hacad184a9;
			11'h370: dataout<=36'h7ddf05cf2;
			11'h371: dataout<=36'h2db3621c2;
			11'h372: dataout<=36'h92b92f56a;
			11'h373: dataout<=36'haa9ed7d74;
			11'h374: dataout<=36'h7dbf05fa1;
			11'h375: dataout<=36'h2ef9623bb;
			11'h376: dataout<=36'h93cd6ee74;
			11'h377: dataout<=36'ha89a97612;
			11'h378: dataout<=36'h7d9dc6251;
			11'h379: dataout<=36'h303e625c4;
			11'h37a: dataout<=36'h94e9ae78d;
			11'h37b: dataout<=36'ha6a056e85;
			11'h37c: dataout<=36'h7d7bc64ff;
			11'h37d: dataout<=36'h3181a27da;
			11'h37e: dataout<=36'h960c6e0ba;
			11'h37f: dataout<=36'ha4b0966ce;
			11'h380: dataout<=36'h7d58c67ad;
			11'h381: dataout<=36'h32c3a29ff;
			11'h382: dataout<=36'h9736ad9fa;
			11'h383: dataout<=36'ha2cb95eec;
			11'h384: dataout<=36'h7d34c6a5a;
			11'h385: dataout<=36'h340422c32;
			11'h386: dataout<=36'h9867ed34d;
			11'h387: dataout<=36'ha0f1556e1;
			11'h388: dataout<=36'h7d1006d06;
			11'h389: dataout<=36'h354322e71;
			11'h38a: dataout<=36'h999f6ccb3;
			11'h38b: dataout<=36'h9f2254eaf;
			11'h38c: dataout<=36'h7cea46fb1;
			11'h38d: dataout<=36'h3680230be;
			11'h38e: dataout<=36'h9addac630;
			11'h38f: dataout<=36'h9d5e94655;
			11'h390: dataout<=36'h7cc3c725c;
			11'h391: dataout<=36'h37bc63318;
			11'h392: dataout<=36'h9c226bfbd;
			11'h393: dataout<=36'h9ba653dd5;
			11'h394: dataout<=36'h7c9c47506;
			11'h395: dataout<=36'h38f6a3580;
			11'h396: dataout<=36'h9d6deb961;
			11'h397: dataout<=36'h99f9d3530;
			11'h398: dataout<=36'h7c73c77ae;
			11'h399: dataout<=36'h3a2ea37f6;
			11'h39a: dataout<=36'h9ebfeb31e;
			11'h39b: dataout<=36'h985912c67;
			11'h39c: dataout<=36'h7c4a87a56;
			11'h39d: dataout<=36'h3b65a3a78;
			11'h39e: dataout<=36'ha0182aced;
			11'h39f: dataout<=36'h96c49237a;
			11'h3a0: dataout<=36'h7c2007cfd;
			11'h3a1: dataout<=36'h3c9a63d0a;
			11'h3a2: dataout<=36'ha1776a6d5;
			11'h3a3: dataout<=36'h953c51a6c;
			11'h3a4: dataout<=36'h7bf507fa4;
			11'h3a5: dataout<=36'h3dce63fa6;
			11'h3a6: dataout<=36'ha2dc2a0ce;
			11'h3a7: dataout<=36'h93c09113d;
			11'h3a8: dataout<=36'h7bc908249;
			11'h3a9: dataout<=36'h3effa4250;
			11'h3aa: dataout<=36'ha44729ae3;
			11'h3ab: dataout<=36'h9251907ee;
			11'h3ac: dataout<=36'h7b9c084ed;
			11'h3ad: dataout<=36'h402f24507;
			11'h3ae: dataout<=36'ha5b7e950f;
			11'h3af: dataout<=36'h90ef0fe80;
			11'h3b0: dataout<=36'h7b6e08791;
			11'h3b1: dataout<=36'h415d247cd;
			11'h3b2: dataout<=36'ha72fa8f52;
			11'h3b3: dataout<=36'h8f99cf4f4;
			11'h3b4: dataout<=36'h7b3f48a33;
			11'h3b5: dataout<=36'h4288e4a9e;
			11'h3b6: dataout<=36'ha8ac689ae;
			11'h3b7: dataout<=36'h8e518eb4c;
			11'h3b8: dataout<=36'h7b0f88cd4;
			11'h3b9: dataout<=36'h43b2a4d7c;
			11'h3ba: dataout<=36'haa2ee8423;
			11'h3bb: dataout<=36'h8d168e188;
			11'h3bc: dataout<=36'h7adf08f75;
			11'h3bd: dataout<=36'h44db25066;
			11'h3be: dataout<=36'habb727ead;
			11'h3bf: dataout<=36'h8be90d7aa;
			11'h3c0: dataout<=36'h7aad89214;
			11'h3c1: dataout<=36'h4600e535e;
			11'h3c2: dataout<=36'had4527955;
			11'h3c3: dataout<=36'h8ac90cdb3;
			11'h3c4: dataout<=36'h7a7b494b2;
			11'h3c5: dataout<=36'h4724a5660;
			11'h3c6: dataout<=36'haed7a7415;
			11'h3c7: dataout<=36'h89b6cc3a4;
			11'h3c8: dataout<=36'h7a480974f;
			11'h3c9: dataout<=36'h4846a5970;
			11'h3ca: dataout<=36'hb07026eee;
			11'h3cb: dataout<=36'h88b24b97e;
			11'h3cc: dataout<=36'h7a13c99eb;
			11'h3cd: dataout<=36'h496625c8e;
			11'h3ce: dataout<=36'hb20e669e4;
			11'h3cf: dataout<=36'h87bbcaf42;
			11'h3d0: dataout<=36'h79dec9c86;
			11'h3d1: dataout<=36'h4a83e5fb6;
			11'h3d2: dataout<=36'hb3b0e64f2;
			11'h3d3: dataout<=36'h86d34a4f2;
			11'h3d4: dataout<=36'h79a8c9f20;
			11'h3d5: dataout<=36'h4b9f662ec;
			11'h3d6: dataout<=36'hb5596601c;
			11'h3d7: dataout<=36'h85f8c9a8e;
			11'h3d8: dataout<=36'h79720a1b8;
			11'h3d9: dataout<=36'h4cb86662c;
			11'h3da: dataout<=36'hb705a5b62;
			11'h3db: dataout<=36'h852cc9019;
			11'h3dc: dataout<=36'h793a4a450;
			11'h3dd: dataout<=36'h4dcfa6979;
			11'h3de: dataout<=36'hb8b7656c1;
			11'h3df: dataout<=36'h846f08593;
			11'h3e0: dataout<=36'h7901ca6e6;
			11'h3e1: dataout<=36'h4ee426cd1;
			11'h3e2: dataout<=36'hba6d6523e;
			11'h3e3: dataout<=36'h83bf87afd;
			11'h3e4: dataout<=36'h78c84a97b;
			11'h3e5: dataout<=36'h4ff6a7036;
			11'h3e6: dataout<=36'hbc2864dd7;
			11'h3e7: dataout<=36'h831ec7058;
			11'h3e8: dataout<=36'h788dcac0f;
			11'h3e9: dataout<=36'h5106a73a7;
			11'h3ea: dataout<=36'hbde7e498d;
			11'h3eb: dataout<=36'h828c865a7;
			11'h3ec: dataout<=36'h78528aea1;
			11'h3ed: dataout<=36'h521427723;
			11'h3ee: dataout<=36'hbfab64561;
			11'h3ef: dataout<=36'h8208c5aea;
			11'h3f0: dataout<=36'h78168b132;
			11'h3f1: dataout<=36'h531f67aa9;
			11'h3f2: dataout<=36'hc172e4150;
			11'h3f3: dataout<=36'h819405022;
			11'h3f4: dataout<=36'h77d98b3c2;
			11'h3f5: dataout<=36'h542827e3c;
			11'h3f6: dataout<=36'hc33ee3d5d;
			11'h3f7: dataout<=36'h812dc4550;
			11'h3f8: dataout<=36'h779bcb651;
			11'h3f9: dataout<=36'h552ee81d9;
			11'h3fa: dataout<=36'hc50ee3985;
			11'h3fb: dataout<=36'h80d683a77;
			11'h3fc: dataout<=36'h775d0b8de;
			11'h3fd: dataout<=36'h5632a8582;
			11'h3fe: dataout<=36'hc6e2635ce;
			11'h3ff: dataout<=36'h808e02f97;
			11'h400: dataout<=36'h771d4bb6a;
			11'h401: dataout<=36'h573428937;
			11'h402: dataout<=36'hc8ba63235;
			11'h403: dataout<=36'h8054824b1;
			11'h404: dataout<=36'h76dccbdf5;
			11'h405: dataout<=36'h583328cf7;
			11'h406: dataout<=36'hca95e2eb9;
			11'h407: dataout<=36'h8029c19c7;
			11'h408: dataout<=36'h769b8c07e;
			11'h409: dataout<=36'h592f690c0;
			11'h40a: dataout<=36'hcc7462b5c;
			11'h40b: dataout<=36'h800e00eda;
			11'h40c: dataout<=36'h76594c306;
			11'h40d: dataout<=36'h5a2929495;
			11'h40e: dataout<=36'hce56a281e;
			11'h40f: dataout<=36'h8001003eb;
			11'h410: dataout<=36'h76164c58c;
			11'h411: dataout<=36'h5b2029873;
			11'h412: dataout<=36'hd03ba24ff;
			11'h413: dataout<=36'h80037f8fd;
			11'h414: dataout<=36'h75d24c811;
			11'h415: dataout<=36'h5c1469c5d;
			11'h416: dataout<=36'hd22422200;
			11'h417: dataout<=36'h80147ee0f;
			11'h418: dataout<=36'h758d8ca94;
			11'h419: dataout<=36'h5d05ea051;
			11'h41a: dataout<=36'hd40f61f20;
			11'h41b: dataout<=36'h80347e322;
			11'h41c: dataout<=36'h7547ccd16;
			11'h41d: dataout<=36'h5df4ea450;
			11'h41e: dataout<=36'hd5fe21c60;
			11'h41f: dataout<=36'h80637d83a;
			11'h420: dataout<=36'h75014cf97;
			11'h421: dataout<=36'h5ee16a859;
			11'h422: dataout<=36'hd7efa19bd;
			11'h423: dataout<=36'h80a13cd55;
			11'h424: dataout<=36'h74ba0d216;
			11'h425: dataout<=36'h5fcaeac6a;
			11'h426: dataout<=36'hd9e2e173b;
			11'h427: dataout<=36'h80edfc277;
			11'h428: dataout<=36'h7471cd493;
			11'h429: dataout<=36'h60b16b087;
			11'h42a: dataout<=36'hdbd9214db;
			11'h42b: dataout<=36'h81497b7a0;
			11'h42c: dataout<=36'h7428cd70f;
			11'h42d: dataout<=36'h61956b4ac;
			11'h42e: dataout<=36'hddd1a1299;
			11'h42f: dataout<=36'h81b3bacd1;
			11'h430: dataout<=36'h73decd989;
			11'h431: dataout<=36'h62762b8dd;
			11'h432: dataout<=36'hdfcca107b;
			11'h433: dataout<=36'h822cba20c;
			11'h434: dataout<=36'h73940dc02;
			11'h435: dataout<=36'h63546bd16;
			11'h436: dataout<=36'he1c9a0e7a;
			11'h437: dataout<=36'h82b479752;
			11'h438: dataout<=36'h73484de79;
			11'h439: dataout<=36'h642f6c15a;
			11'h43a: dataout<=36'he3c8e0c9d;
			11'h43b: dataout<=36'h834af8ca4;
			11'h43c: dataout<=36'h72fc0e0ef;
			11'h43d: dataout<=36'h65082c5a5;
			11'h43e: dataout<=36'he5c9a0adb;
			11'h43f: dataout<=36'h83eff8204;
			11'h440: dataout<=36'h72aece362;
			11'h441: dataout<=36'h65dd2c9fa;
			11'h442: dataout<=36'he7cbe0940;
			11'h443: dataout<=36'h84a337772;
			11'h444: dataout<=36'h72608e5d5;
			11'h445: dataout<=36'h66afece5a;
			11'h446: dataout<=36'he9d0e07c2;
			11'h447: dataout<=36'h856536cf0;
			11'h448: dataout<=36'h72118e845;
			11'h449: dataout<=36'h677eed2c1;
			11'h44a: dataout<=36'hebd620669;
			11'h44b: dataout<=36'h863536280;
			11'h44c: dataout<=36'h71c1ceab4;
			11'h44d: dataout<=36'h684b6d731;
			11'h44e: dataout<=36'heddd2052e;
			11'h44f: dataout<=36'h8713b5822;
			11'h450: dataout<=36'h71714ed21;
			11'h451: dataout<=36'h6914edba9;
			11'h452: dataout<=36'hefe520414;
			11'h453: dataout<=36'h880034dd7;
			11'h454: dataout<=36'h711fcef8c;
			11'h455: dataout<=36'h69daee02a;
			11'h456: dataout<=36'hf1ee2031e;
			11'h457: dataout<=36'h88fab43a1;
			11'h458: dataout<=36'h70cd8f1f6;
			11'h459: dataout<=36'h6a9e2e4b4;
			11'h45a: dataout<=36'hf3f860247;
			11'h45b: dataout<=36'h8a0333982;
			11'h45c: dataout<=36'h707a4f45e;
			11'h45d: dataout<=36'h6b5e2e947;
			11'h45e: dataout<=36'hf603a0194;
			11'h45f: dataout<=36'h8b1932f79;
			11'h460: dataout<=36'h70268f6c4;
			11'h461: dataout<=36'h6c1b2ede0;
			11'h462: dataout<=36'hf80ee00ff;
			11'h463: dataout<=36'h8c3d32589;
			11'h464: dataout<=36'h6fd1cf928;
			11'h465: dataout<=36'h6cd4ef282;
			11'h466: dataout<=36'hfa1ae008e;
			11'h467: dataout<=36'h8d6e71bb2;
			11'h468: dataout<=36'h6f7c4fb8b;
			11'h469: dataout<=36'h6d8baf72c;
			11'h46a: dataout<=36'hfc276003d;
			11'h46b: dataout<=36'h8ead311f6;
			11'h46c: dataout<=36'h6f25cfdeb;
			11'h46d: dataout<=36'h6e3eafbde;
			11'h46e: dataout<=36'hfe3420011;
			11'h46f: dataout<=36'h8ff930856;
			11'h470: dataout<=36'h6eced004a;
			11'h471: dataout<=36'h6eef30097;
			11'h472: dataout<=36'h0040e0002;
			11'h473: dataout<=36'h91522fed2;
			11'h474: dataout<=36'h6e76d02a7;
			11'h475: dataout<=36'h6f9c30558;
			11'h476: dataout<=36'h024de0017;
			11'h477: dataout<=36'h92b82f56d;
			11'h478: dataout<=36'h6e1dd0502;
			11'h479: dataout<=36'h7045b0a21;
			11'h47a: dataout<=36'h045ae0050;
			11'h47b: dataout<=36'h942aeec27;
			11'h47c: dataout<=36'h6dc45075b;
			11'h47d: dataout<=36'h70ebf0ef0;
			11'h47e: dataout<=36'h0666e00a8;
			11'h47f: dataout<=36'h95aa2e301;
			11'h480: dataout<=36'h6d69d09b2;
			11'h481: dataout<=36'h718ef13c6;
			11'h482: dataout<=36'h0872e0122;
			11'h483: dataout<=36'h9735ed9fc;
			11'h484: dataout<=36'h6d0ed0c07;
			11'h485: dataout<=36'h722ef18a2;
			11'h486: dataout<=36'h0a7de01bc;
			11'h487: dataout<=36'h98cded11a;
			11'h488: dataout<=36'h6cb2d0e5b;
			11'h489: dataout<=36'h72cbb1d87;
			11'h48a: dataout<=36'h0c8920278;
			11'h48b: dataout<=36'h9a71ec85b;
			11'h48c: dataout<=36'h6c56110ac;
			11'h48d: dataout<=36'h7364b2271;
			11'h48e: dataout<=36'h0e92e0356;
			11'h48f: dataout<=36'h9c21abfc0;
			11'h490: dataout<=36'h6bf8512fb;
			11'h491: dataout<=36'h73f9f2763;
			11'h492: dataout<=36'h109be0459;
			11'h493: dataout<=36'h9ddd2b74b;
			11'h494: dataout<=36'h6b9a11549;
			11'h495: dataout<=36'h748cb2c5a;
			11'h496: dataout<=36'h12a3e0578;
			11'h497: dataout<=36'h9fa42aefc;
			11'h498: dataout<=36'h6b3ad1794;
			11'h499: dataout<=36'h751b73158;
			11'h49a: dataout<=36'h14aaa06bc;
			11'h49b: dataout<=36'ha1766a6d5;
			11'h49c: dataout<=36'h6adb119dd;
			11'h49d: dataout<=36'h75a6f365a;
			11'h49e: dataout<=36'h16af6081e;
			11'h49f: dataout<=36'ha353a9ed5;
			11'h4a0: dataout<=36'h6a7a51c24;
			11'h4a1: dataout<=36'h762ef3b63;
			11'h4a2: dataout<=36'h18b2e09a3;
			11'h4a3: dataout<=36'ha53be96ff;
			11'h4a4: dataout<=36'h6a18d1e6a;
			11'h4a5: dataout<=36'h76b3f4074;
			11'h4a6: dataout<=36'h1ab5e0b48;
			11'h4a7: dataout<=36'ha72e68f54;
			11'h4a8: dataout<=36'h69b6920ad;
			11'h4a9: dataout<=36'h773534588;
			11'h4aa: dataout<=36'h1cb620d0e;
			11'h4ab: dataout<=36'ha92ba87d3;
			11'h4ac: dataout<=36'h6953922ee;
			11'h4ad: dataout<=36'h77b2f4aa2;
			11'h4ae: dataout<=36'h1eb4a0ef5;
			11'h4af: dataout<=36'hab32a807e;
			11'h4b0: dataout<=36'h68efd252c;
			11'h4b1: dataout<=36'h782cf4fc1;
			11'h4b2: dataout<=36'h20b0e10fd;
			11'h4b3: dataout<=36'had43e7956;
			11'h4b4: dataout<=36'h688b12769;
			11'h4b5: dataout<=36'h78a3754e7;
			11'h4b6: dataout<=36'h22ab61328;
			11'h4b7: dataout<=36'haf5ea725b;
			11'h4b8: dataout<=36'h6825d29a3;
			11'h4b9: dataout<=36'h791675a10;
			11'h4ba: dataout<=36'h24a321571;
			11'h4bb: dataout<=36'hb182e6b8f;
			11'h4bc: dataout<=36'h67bfd2bdc;
			11'h4bd: dataout<=36'h798675f3e;
			11'h4be: dataout<=36'h2699217d8;
			11'h4bf: dataout<=36'hb3b0264f3;
			11'h4c0: dataout<=36'h6758d2e12;
			11'h4c1: dataout<=36'h79f276472;
			11'h4c2: dataout<=36'h288c61a62;
			11'h4c3: dataout<=36'hb5e665e86;
			11'h4c4: dataout<=36'h66f153046;
			11'h4c5: dataout<=36'h7a5af69a9;
			11'h4c6: dataout<=36'h2a7ca1d0a;
			11'h4c7: dataout<=36'hb8256584a;
			11'h4c8: dataout<=36'h6688d3278;
			11'h4c9: dataout<=36'h7abff6ee7;
			11'h4ca: dataout<=36'h2c6ae1fd5;
			11'h4cb: dataout<=36'hba6ca523f;
			11'h4cc: dataout<=36'h661fd34a7;
			11'h4cd: dataout<=36'h7b2137426;
			11'h4ce: dataout<=36'h2e55222bc;
			11'h4cf: dataout<=36'hbcbc24c67;
			11'h4d0: dataout<=36'h65b6136d4;
			11'h4d1: dataout<=36'h7b7ef7969;
			11'h4d2: dataout<=36'h303c625c3;
			11'h4d3: dataout<=36'hbf13646c1;
			11'h4d4: dataout<=36'h654b538ff;
			11'h4d5: dataout<=36'h7bd8f7eb3;
			11'h4d6: dataout<=36'h3221228ec;
			11'h4d7: dataout<=36'hc1722414f;
			11'h4d8: dataout<=36'h64e013b28;
			11'h4d9: dataout<=36'h7c2fb83ff;
			11'h4da: dataout<=36'h3402a2c30;
			11'h4db: dataout<=36'hc3d863c11;
			11'h4dc: dataout<=36'h647413d4e;
			11'h4dd: dataout<=36'h7c82b894e;
			11'h4de: dataout<=36'h35e062f94;
			11'h4df: dataout<=36'hc645a3708;
			11'h4e0: dataout<=36'h640753f72;
			11'h4e1: dataout<=36'h7cd1f8ea1;
			11'h4e2: dataout<=36'h37baa3317;
			11'h4e3: dataout<=36'hc8b963235;
			11'h4e4: dataout<=36'h639994194;
			11'h4e5: dataout<=36'h7d1d793f9;
			11'h4e6: dataout<=36'h3991636ba;
			11'h4e7: dataout<=36'hcb33e2d97;
			11'h4e8: dataout<=36'h632b543b3;
			11'h4e9: dataout<=36'h7d6579952;
			11'h4ea: dataout<=36'h3b6423a79;
			11'h4eb: dataout<=36'hcdb46292f;
			11'h4ec: dataout<=36'h62bc945d1;
			11'h4ed: dataout<=36'h7daa79eaf;
			11'h4ee: dataout<=36'h3d33a3e53;
			11'h4ef: dataout<=36'hd03ae24ff;
			11'h4f0: dataout<=36'h624cd47eb;
			11'h4f1: dataout<=36'h7deaba40e;
			11'h4f2: dataout<=36'h3efe2424f;
			11'h4f3: dataout<=36'hd2c6e2106;
			11'h4f4: dataout<=36'h61dc54a03;
			11'h4f5: dataout<=36'h7e277a970;
			11'h4f6: dataout<=36'h40c4a4668;
			11'h4f7: dataout<=36'hd55821d45;
			11'h4f8: dataout<=36'h616b54c19;
			11'h4f9: dataout<=36'h7e60faed4;
			11'h4fa: dataout<=36'h428764a9b;
			11'h4fb: dataout<=36'hd7ee619bd;
			11'h4fc: dataout<=36'h60f954e2d;
			11'h4fd: dataout<=36'h7e96bb43d;
			11'h4fe: dataout<=36'h444624eee;
			11'h4ff: dataout<=36'hda896166d;
			11'h500: dataout<=36'h6086d503e;
			11'h501: dataout<=36'h7ec8bb9a6;
			11'h502: dataout<=36'h45ffe535b;
			11'h503: dataout<=36'hdd28a1356;
			11'h504: dataout<=36'h60139524c;
			11'h505: dataout<=36'h7ef6bbf11;
			11'h506: dataout<=36'h47b4a57e6;
			11'h507: dataout<=36'hdfcbe1079;
			11'h508: dataout<=36'h5f9f95458;
			11'h509: dataout<=36'h7f213c47e;
			11'h50a: dataout<=36'h4964e5c8c;
			11'h50b: dataout<=36'he27320dd5;
			11'h50c: dataout<=36'h5f2b15662;
			11'h50d: dataout<=36'h7f483c9ed;
			11'h50e: dataout<=36'h4b10a614d;
			11'h50f: dataout<=36'he51da0b6c;
			11'h510: dataout<=36'h5eb595869;
			11'h511: dataout<=36'h7f6b3cf5e;
			11'h512: dataout<=36'h4cb76662b;
			11'h513: dataout<=36'he7cb6093e;
			11'h514: dataout<=36'h5e3f95a6d;
			11'h515: dataout<=36'h7f8a7d4cf;
			11'h516: dataout<=36'h4e5866b22;
			11'h517: dataout<=36'hea7be074a;
			11'h518: dataout<=36'h5dc8d5c6f;
			11'h519: dataout<=36'h7fa5fda43;
			11'h51a: dataout<=36'h4ff4e7035;
			11'h51b: dataout<=36'hed2f20591;
			11'h51c: dataout<=36'h5d5195e6f;
			11'h51d: dataout<=36'h7fbe3dfb7;
			11'h51e: dataout<=36'h518c67560;
			11'h51f: dataout<=36'hefe460413;
			11'h520: dataout<=36'h5cd95606c;
			11'h521: dataout<=36'h7fd23e52d;
			11'h522: dataout<=36'h531e67aa8;
			11'h523: dataout<=36'hf29b602d0;
			11'h524: dataout<=36'h5c6096266;
			11'h525: dataout<=36'h7fe2beaa3;
			11'h526: dataout<=36'h54aaa8008;
			11'h527: dataout<=36'hf554201c9;
			11'h528: dataout<=36'h5be71645e;
			11'h529: dataout<=36'h7fef7f01a;
			11'h52a: dataout<=36'h5631a8582;
			11'h52b: dataout<=36'hf80e200fd;
			11'h52c: dataout<=36'h5b6d16653;
			11'h52d: dataout<=36'h7ff87f590;
			11'h52e: dataout<=36'h57b268b13;
			11'h52f: dataout<=36'hfac8e006d;
			11'h530: dataout<=36'h5af256846;
			11'h531: dataout<=36'h7ffdffb08;
			11'h532: dataout<=36'h592e290bd;
			11'h533: dataout<=36'hfd8460019;
			11'h534: dataout<=36'h5a76d6a36;
			11'h535: dataout<=36'h7fff40080;
			11'h536: dataout<=36'h5aa3e9680;
			11'h537: dataout<=36'h004020001;
			11'h538: dataout<=36'h59fad6c23;
			11'h539: dataout<=36'h7ffd005f7;
			11'h53a: dataout<=36'h5c1329c5a;
			11'h53b: dataout<=36'h02fbe0024;
			11'h53c: dataout<=36'h597e16e0e;
			11'h53d: dataout<=36'h7ff740b6f;
			11'h53e: dataout<=36'h5d7d2a24c;
			11'h53f: dataout<=36'h05b720083;
			11'h540: dataout<=36'h590096ff6;
			11'h541: dataout<=36'h7fed810e6;
			11'h542: dataout<=36'h5ee06a855;
			11'h543: dataout<=36'h0871e011e;
			11'h544: dataout<=36'h5882971db;
			11'h545: dataout<=36'h7fe00165c;
			11'h546: dataout<=36'h603d6ae74;
			11'h547: dataout<=36'h0b2ba01f5;
			11'h548: dataout<=36'h5803d73bd;
			11'h549: dataout<=36'h7fcec1bd2;
			11'h54a: dataout<=36'h61942b4aa;
			11'h54b: dataout<=36'h0de420307;
			11'h54c: dataout<=36'h57849759d;
			11'h54d: dataout<=36'h7fba02146;
			11'h54e: dataout<=36'h62e46baf4;
			11'h54f: dataout<=36'h109ae0454;
			11'h550: dataout<=36'h57049777a;
			11'h551: dataout<=36'h7fa1426ba;
			11'h552: dataout<=36'h642e2c155;
			11'h553: dataout<=36'h134fe05dd;
			11'h554: dataout<=36'h5683d7955;
			11'h555: dataout<=36'h7f8502c2f;
			11'h556: dataout<=36'h65722c7cc;
			11'h557: dataout<=36'h1602607a1;
			11'h558: dataout<=36'h560297b2c;
			11'h559: dataout<=36'h7f64c31a0;
			11'h55a: dataout<=36'h66ae6ce56;
			11'h55b: dataout<=36'h18b26099f;
			11'h55c: dataout<=36'h5580d7d01;
			11'h55d: dataout<=36'h7f4143710;
			11'h55e: dataout<=36'h67e4ad4f3;
			11'h55f: dataout<=36'h1b5fa0bd9;
			11'h560: dataout<=36'h54fe57ed3;
			11'h561: dataout<=36'h7f19c3c7e;
			11'h562: dataout<=36'h6913adba4;
			11'h563: dataout<=36'h1e09a0e4d;
			11'h564: dataout<=36'h547b180a3;
			11'h565: dataout<=36'h7eee841ed;
			11'h566: dataout<=36'h6a3c6e26b;
			11'h567: dataout<=36'h20b0210fb;
			11'h568: dataout<=36'h53f75826f;
			11'h569: dataout<=36'h7ebf84757;
			11'h56a: dataout<=36'h6b5d2e943;
			11'h56b: dataout<=36'h2352e13e2;
			11'h56c: dataout<=36'h537318439;
			11'h56d: dataout<=36'h7e8d04cc0;
			11'h56e: dataout<=36'h6c77af02c;
			11'h56f: dataout<=36'h25f161703;
			11'h570: dataout<=36'h52ee18600;
			11'h571: dataout<=36'h7e56c5227;
			11'h572: dataout<=36'h6d8aef728;
			11'h573: dataout<=36'h288b61a5e;
			11'h574: dataout<=36'h5268587c4;
			11'h575: dataout<=36'h7e1c8578c;
			11'h576: dataout<=36'h6e96afe38;
			11'h577: dataout<=36'h2b20e1df1;
			11'h578: dataout<=36'h51e258985;
			11'h579: dataout<=36'h7ddf05ced;
			11'h57a: dataout<=36'h6f9b30554;
			11'h57b: dataout<=36'h2db1221bc;
			11'h57c: dataout<=36'h515b98b43;
			11'h57d: dataout<=36'h7d9dc624b;
			11'h57e: dataout<=36'h709870c82;
			11'h57f: dataout<=36'h303c225bf;
			11'h580: dataout<=36'h50d418cfe;
			11'h581: dataout<=36'h7d58467a8;
			11'h582: dataout<=36'h718df13c3;
			11'h583: dataout<=36'h32c1629fa;
			11'h584: dataout<=36'h504c18eb7;
			11'h585: dataout<=36'h7d0fc6d02;
			11'h586: dataout<=36'h727cb1b12;
			11'h587: dataout<=36'h3540e2e6b;
			11'h588: dataout<=36'h4fc39906c;
			11'h589: dataout<=36'h7cc347257;
			11'h58a: dataout<=36'h73633226f;
			11'h58b: dataout<=36'h37ba23313;
			11'h58c: dataout<=36'h4f3a9921f;
			11'h58d: dataout<=36'h7c73c77a9;
			11'h58e: dataout<=36'h7442f29d8;
			11'h58f: dataout<=36'h3a2ce37f0;
			11'h590: dataout<=36'h4eb0d93cf;
			11'h591: dataout<=36'h7c2007cf9;
			11'h592: dataout<=36'h751af3154;
			11'h593: dataout<=36'h3c98e3d03;
			11'h594: dataout<=36'h4e269957b;
			11'h595: dataout<=36'h7bc8c8243;
			11'h596: dataout<=36'h75ea738da;
			11'h597: dataout<=36'h3efda424a;
			11'h598: dataout<=36'h4d9bd9725;
			11'h599: dataout<=36'h7b6e0878b;
			11'h59a: dataout<=36'h76b2f406e;
			11'h59b: dataout<=36'h415b247c6;
			11'h59c: dataout<=36'h4d10598cc;
			11'h59d: dataout<=36'h7b0f88ccf;
			11'h59e: dataout<=36'h777374810;
			11'h59f: dataout<=36'h43b0e4d75;
			11'h5a0: dataout<=36'h4c8459a70;
			11'h5a1: dataout<=36'h7aad8920f;
			11'h5a2: dataout<=36'h782c34fbe;
			11'h5a3: dataout<=36'h45fee5356;
			11'h5a4: dataout<=36'h4bf7d9c11;
			11'h5a5: dataout<=36'h7a480974a;
			11'h5a6: dataout<=36'h78dcf5776;
			11'h5a7: dataout<=36'h4844a596a;
			11'h5a8: dataout<=36'h4b6ad9daf;
			11'h5a9: dataout<=36'h79df09c81;
			11'h5aa: dataout<=36'h7985f5f39;
			11'h5ab: dataout<=36'h4a8225faf;
			11'h5ac: dataout<=36'h4add19f4a;
			11'h5ad: dataout<=36'h79724a1b4;
			11'h5ae: dataout<=36'h7a26f6709;
			11'h5af: dataout<=36'h4cb6a6625;
			11'h5b0: dataout<=36'h4a4eda0e1;
			11'h5b1: dataout<=36'h79018a6e1;
			11'h5b2: dataout<=36'h7abef6ee2;
			11'h5b3: dataout<=36'h4ee266cca;
			11'h5b4: dataout<=36'h49c01a276;
			11'h5b5: dataout<=36'h788dcac0a;
			11'h5b6: dataout<=36'h7b4ff76c4;
			11'h5b7: dataout<=36'h5104e739f;
			11'h5b8: dataout<=36'h4930da408;
			11'h5b9: dataout<=36'h78168b12e;
			11'h5ba: dataout<=36'h7bd8b7eaf;
			11'h5bb: dataout<=36'h531de7aa2;
			11'h5bc: dataout<=36'h48a11a596;
			11'h5bd: dataout<=36'h779b8b64b;
			11'h5be: dataout<=36'h7c58b86a1;
			11'h5bf: dataout<=36'h552d281d2;
			11'h5c0: dataout<=36'h4810da722;
			11'h5c1: dataout<=36'h771d8bb65;
			11'h5c2: dataout<=36'h7cd178e9d;
			11'h5c3: dataout<=36'h5732a892f;
			11'h5c4: dataout<=36'h477fda8aa;
			11'h5c5: dataout<=36'h769b4c079;
			11'h5c6: dataout<=36'h7d41396a1;
			11'h5c7: dataout<=36'h592de90b8;
			11'h5c8: dataout<=36'h46ee9aa30;
			11'h5c9: dataout<=36'h76168c587;
			11'h5ca: dataout<=36'h7da9b9ea9;
			11'h5cb: dataout<=36'h5b1ea986b;
			11'h5cc: dataout<=36'h465c9abb2;
			11'h5cd: dataout<=36'h758d8ca90;
			11'h5ce: dataout<=36'h7e08fa6bb;
			11'h5cf: dataout<=36'h5d04aa049;
			11'h5d0: dataout<=36'h45ca5ad31;
			11'h5d1: dataout<=36'h75018cf91;
			11'h5d2: dataout<=36'h7e607aecf;
			11'h5d3: dataout<=36'h5edfea84f;
			11'h5d4: dataout<=36'h45375aead;
			11'h5d5: dataout<=36'h7471cd48e;
			11'h5d6: dataout<=36'h7eaf7b6ec;
			11'h5d7: dataout<=36'h60b02b07e;
			11'h5d8: dataout<=36'h44a3db026;
			11'h5d9: dataout<=36'h73decd985;
			11'h5da: dataout<=36'h7ef63bf0d;
			11'h5db: dataout<=36'h62752b8d4;
			11'h5dc: dataout<=36'h44101b19c;
			11'h5dd: dataout<=36'h7348cde74;
			11'h5de: dataout<=36'h7f34fc730;
			11'h5df: dataout<=36'h642e6c150;
			11'h5e0: dataout<=36'h437b9b30e;
			11'h5e1: dataout<=36'h72aece35d;
			11'h5e2: dataout<=36'h7f6a7cf58;
			11'h5e3: dataout<=36'h65dc2c9f2;
			11'h5e4: dataout<=36'h42e69b47e;
			11'h5e5: dataout<=36'h7211ce841;
			11'h5e6: dataout<=36'h7f987d785;
			11'h5e7: dataout<=36'h677e2d2b7;
			11'h5e8: dataout<=36'h42515b5ea;
			11'h5e9: dataout<=36'h71718ed1c;
			11'h5ea: dataout<=36'h7fbdfdfb2;
			11'h5eb: dataout<=36'h6913edba0;
			11'h5ec: dataout<=36'h41bb5b753;
			11'h5ed: dataout<=36'h70cdcf1f2;
			11'h5ee: dataout<=36'h7fdabe7e3;
			11'h5ef: dataout<=36'h6a9d2e4ab;
			11'h5f0: dataout<=36'h41251b8b9;
			11'h5f1: dataout<=36'h70270f6c0;
			11'h5f2: dataout<=36'h7fefbf014;
			11'h5f3: dataout<=36'h6c1a2edd7;
			11'h5f4: dataout<=36'h408e1ba1b;
			11'h5f5: dataout<=36'h6f7c4fb86;
			11'h5f6: dataout<=36'h7ffaff848;
			11'h5f7: dataout<=36'h6d8aaf723;
			11'h5f8: dataout<=36'h3ff6dbb7b;
			11'h5f9: dataout<=36'h6ecf10046;
			11'h5fa: dataout<=36'h7fff0007b;
			11'h5fb: dataout<=36'h6eee7008e;
			11'h5fc: dataout<=36'h3f5f1bcd7;
			11'h5fd: dataout<=36'h6e1e504fe;
			11'h5fe: dataout<=36'h7ffa408af;
			11'h5ff: dataout<=36'h7044f0a16;
			11'h600: dataout<=36'h3ec6dbe2f;
			11'h601: dataout<=36'h6d6a109ad;
			11'h602: dataout<=36'h7fecc10e0;
			11'h603: dataout<=36'h718e713bc;
			11'h604: dataout<=36'h3e2e1bf85;
			11'h605: dataout<=36'h6cb2d0e56;
			11'h606: dataout<=36'h7fd741913;
			11'h607: dataout<=36'h72cab1d7d;
			11'h608: dataout<=36'h3d951c0d7;
			11'h609: dataout<=36'h6bf8d12f6;
			11'h60a: dataout<=36'h7fb982141;
			11'h60b: dataout<=36'h73f9b2758;
			11'h60c: dataout<=36'h3cfb5c226;
			11'h60d: dataout<=36'h6b3b1178f;
			11'h60e: dataout<=36'h7f9302970;
			11'h60f: dataout<=36'h751af314d;
			11'h610: dataout<=36'h3c615c372;
			11'h611: dataout<=36'h6a7a91c20;
			11'h612: dataout<=36'h7f648319b;
			11'h613: dataout<=36'h762eb3b5a;
			11'h614: dataout<=36'h3bc6dc4bb;
			11'h615: dataout<=36'h69b6d20a9;
			11'h616: dataout<=36'h7f2dc39c4;
			11'h617: dataout<=36'h7734b457e;
			11'h618: dataout<=36'h3b2c1c600;
			11'h619: dataout<=36'h68f052527;
			11'h61a: dataout<=36'h7eee841e6;
			11'h61b: dataout<=36'h782c74fb7;
			11'h61c: dataout<=36'h3a909c742;
			11'h61d: dataout<=36'h68265299f;
			11'h61e: dataout<=36'h7ea6c4a07;
			11'h61f: dataout<=36'h791675a06;
			11'h620: dataout<=36'h39f4dc880;
			11'h621: dataout<=36'h675952e0d;
			11'h622: dataout<=36'h7e5685221;
			11'h623: dataout<=36'h79f236467;
			11'h624: dataout<=36'h39589c9bc;
			11'h625: dataout<=36'h668953274;
			11'h626: dataout<=36'h7dfe45a38;
			11'h627: dataout<=36'h7abfb6edb;
			11'h628: dataout<=36'h38bc1caf3;
			11'h629: dataout<=36'h65b6936cf;
			11'h62a: dataout<=36'h7d9d86245;
			11'h62b: dataout<=36'h7b7ef7960;
			11'h62c: dataout<=36'h381f1cc28;
			11'h62d: dataout<=36'h64e0d3b23;
			11'h62e: dataout<=36'h7d3506a4e;
			11'h62f: dataout<=36'h7c2fb83f4;
			11'h630: dataout<=36'h37819cd59;
			11'h631: dataout<=36'h6407d3f6e;
			11'h632: dataout<=36'h7cc3c7251;
			11'h633: dataout<=36'h7cd1f8e97;
			11'h634: dataout<=36'h36e39ce87;
			11'h635: dataout<=36'h632bd43b0;
			11'h636: dataout<=36'h7c4a47a4e;
			11'h637: dataout<=36'h7d65b9947;
			11'h638: dataout<=36'h36455cfb1;
			11'h639: dataout<=36'h624d147e7;
			11'h63a: dataout<=36'h7bc88823f;
			11'h63b: dataout<=36'h7deafa403;
			11'h63c: dataout<=36'h35a6dd0d8;
			11'h63d: dataout<=36'h616bd4c14;
			11'h63e: dataout<=36'h7b3f48a27;
			11'h63f: dataout<=36'h7e613aeca;
			11'h640: dataout<=36'h3507dd1fc;
			11'h641: dataout<=36'h608795039;
			11'h642: dataout<=36'h7aadc9209;
			11'h643: dataout<=36'h7ec8fb99b;
			11'h644: dataout<=36'h34685d31c;
			11'h645: dataout<=36'h5fa015453;
			11'h646: dataout<=36'h7a13899e0;
			11'h647: dataout<=36'h7f21bc473;
			11'h648: dataout<=36'h33c89d439;
			11'h649: dataout<=36'h5eb655864;
			11'h64a: dataout<=36'h79724a1ad;
			11'h64b: dataout<=36'h7f6bbcf53;
			11'h64c: dataout<=36'h33285d552;
			11'h64d: dataout<=36'h5dc955c6a;
			11'h64e: dataout<=36'h78c80a970;
			11'h64f: dataout<=36'h7fa6bda38;
			11'h650: dataout<=36'h3287dd668;
			11'h651: dataout<=36'h5cda16067;
			11'h652: dataout<=36'h7816cb127;
			11'h653: dataout<=36'h7fd2fe522;
			11'h654: dataout<=36'h31e6dd77b;
			11'h655: dataout<=36'h5be7d645a;
			11'h656: dataout<=36'h775d4b8d4;
			11'h657: dataout<=36'h7ff03f00e;
			11'h658: dataout<=36'h31459d88a;
			11'h659: dataout<=36'h5af316841;
			11'h65a: dataout<=36'h769c0c073;
			11'h65b: dataout<=36'h7ffe7fafd;
			11'h65c: dataout<=36'h30a3dd996;
			11'h65d: dataout<=36'h59fb56c1f;
			11'h65e: dataout<=36'h75d28c807;
			11'h65f: dataout<=36'h7ffdc05eb;
			11'h660: dataout<=36'h3001dda9e;
			11'h661: dataout<=36'h590116ff2;
			11'h662: dataout<=36'h75018cf8e;
			11'h663: dataout<=36'h7fee010da;
			11'h664: dataout<=36'h2f5f9dba3;
			11'h665: dataout<=36'h5804973ba;
			11'h666: dataout<=36'h74294d706;
			11'h667: dataout<=36'h7fcf81bc6;
			11'h668: dataout<=36'h2ebcddca4;
			11'h669: dataout<=36'h570517776;
			11'h66a: dataout<=36'h7348cde6f;
			11'h66b: dataout<=36'h7fa2426b0;
			11'h66c: dataout<=36'h2e19ddda2;
			11'h66d: dataout<=36'h560357b29;
			11'h66e: dataout<=36'h72614e5cb;
			11'h66f: dataout<=36'h7f65c3195;
			11'h670: dataout<=36'h2d765de9c;
			11'h671: dataout<=36'h54fed7ecf;
			11'h672: dataout<=36'h71718ed17;
			11'h673: dataout<=36'h7f1ac3c74;
			11'h674: dataout<=36'h2cd29df93;
			11'h675: dataout<=36'h53f7d826c;
			11'h676: dataout<=36'h707acf456;
			11'h677: dataout<=36'h7ec08474c;
			11'h678: dataout<=36'h2c2e9e086;
			11'h679: dataout<=36'h52ee985fb;
			11'h67a: dataout<=36'h6f7c8fb81;
			11'h67b: dataout<=36'h7e57c521b;
			11'h67c: dataout<=36'h2b8a5e176;
			11'h67d: dataout<=36'h51e318981;
			11'h67e: dataout<=36'h6e779029d;
			11'h67f: dataout<=36'h7de045ce1;
			11'h680: dataout<=36'h2ae59e262;
			11'h681: dataout<=36'h50d4d8cfa;
			11'h682: dataout<=36'h6d6a909a8;
			11'h683: dataout<=36'h7d5a0679d;
			11'h684: dataout<=36'h2a409e34b;
			11'h685: dataout<=36'h4fc459068;
			11'h686: dataout<=36'h6c56910a2;
			11'h687: dataout<=36'h7cc50724c;
			11'h688: dataout<=36'h299b5e430;
			11'h689: dataout<=36'h4eb1993ca;
			11'h68a: dataout<=36'h6b3b91789;
			11'h68b: dataout<=36'h7c2187ced;
			11'h68c: dataout<=36'h28f59e512;
			11'h68d: dataout<=36'h4d9c59722;
			11'h68e: dataout<=36'h6a1951e61;
			11'h68f: dataout<=36'h7b6f88781;
			11'h690: dataout<=36'h284fde5f0;
			11'h691: dataout<=36'h4c8519a6c;
			11'h692: dataout<=36'h68f092522;
			11'h693: dataout<=36'h7aaf09204;
			11'h694: dataout<=36'h27a99e6cb;
			11'h695: dataout<=36'h4b6b99dab;
			11'h696: dataout<=36'h67c0d2bd3;
			11'h697: dataout<=36'h79e049c76;
			11'h698: dataout<=36'h27031e7a2;
			11'h699: dataout<=36'h4a4f9a0de;
			11'h69a: dataout<=36'h6689d326f;
			11'h69b: dataout<=36'h79034a6d6;
			11'h69c: dataout<=36'h265c5e875;
			11'h69d: dataout<=36'h49319a403;
			11'h69e: dataout<=36'h654c138f5;
			11'h69f: dataout<=36'h78184b123;
			11'h6a0: dataout<=36'h25b55e945;
			11'h6a1: dataout<=36'h48119a71d;
			11'h6a2: dataout<=36'h640813f68;
			11'h6a3: dataout<=36'h771f4bb5b;
			11'h6a4: dataout<=36'h250e1ea12;
			11'h6a5: dataout<=36'h46ef9aa2c;
			11'h6a6: dataout<=36'h62bdd45c7;
			11'h6a7: dataout<=36'h76184c57d;
			11'h6a8: dataout<=36'h24665eadb;
			11'h6a9: dataout<=36'h45cb1ad2e;
			11'h6aa: dataout<=36'h616c54c11;
			11'h6ab: dataout<=36'h75034cf88;
			11'h6ac: dataout<=36'h23be9eba0;
			11'h6ad: dataout<=36'h44a51b023;
			11'h6ae: dataout<=36'h601515243;
			11'h6af: dataout<=36'h73e0cd97a;
			11'h6b0: dataout<=36'h23165ec62;
			11'h6b1: dataout<=36'h437c9b30c;
			11'h6b2: dataout<=36'h5eb715862;
			11'h6b3: dataout<=36'h72b0ce354;
			11'h6b4: dataout<=36'h226e1ed20;
			11'h6b5: dataout<=36'h42525b5e7;
			11'h6b6: dataout<=36'h5d5315e67;
			11'h6b7: dataout<=36'h71738ed12;
			11'h6b8: dataout<=36'h21c55edda;
			11'h6b9: dataout<=36'h4125db8b5;
			11'h6ba: dataout<=36'h5be856455;
			11'h6bb: dataout<=36'h7028cf6b6;
			11'h6bc: dataout<=36'h211c9ee91;
			11'h6bd: dataout<=36'h3ff81bb77;
			11'h6be: dataout<=36'h5a7896a2d;
			11'h6bf: dataout<=36'h6ed11003c;
			11'h6c0: dataout<=36'h20735ef44;
			11'h6c1: dataout<=36'h3ec7dbe2c;
			11'h6c2: dataout<=36'h5901d6fed;
			11'h6c3: dataout<=36'h6d6c909a4;
			11'h6c4: dataout<=36'h1fca1eff4;
			11'h6c5: dataout<=36'h3d961c0d5;
			11'h6c6: dataout<=36'h578617596;
			11'h6c7: dataout<=36'h6bfb112ee;
			11'h6c8: dataout<=36'h1f205f0a0;
			11'h6c9: dataout<=36'h3c621c370;
			11'h6ca: dataout<=36'h5603d7b26;
			11'h6cb: dataout<=36'h6a7d11c17;
			11'h6cc: dataout<=36'h1e769f148;
			11'h6cd: dataout<=36'h3b2cdc5fd;
			11'h6ce: dataout<=36'h547c5809b;
			11'h6cf: dataout<=36'h68f29251f;
			11'h6d0: dataout<=36'h1dcc9f1ed;
			11'h6d1: dataout<=36'h39f5dc87e;
			11'h6d2: dataout<=36'h52ef985f8;
			11'h6d3: dataout<=36'h675bd2e05;
			11'h6d4: dataout<=36'h1d225f28e;
			11'h6d5: dataout<=36'h38bd1caf0;
			11'h6d6: dataout<=36'h515d18b3b;
			11'h6d7: dataout<=36'h65b8d36c7;
			11'h6d8: dataout<=36'h1c77df32b;
			11'h6d9: dataout<=36'h37825cd55;
			11'h6da: dataout<=36'h4fc4d9063;
			11'h6db: dataout<=36'h640a53f66;
			11'h6dc: dataout<=36'h1bcd1f3c5;
			11'h6dd: dataout<=36'h36465cfae;
			11'h6de: dataout<=36'h4e2819574;
			11'h6df: dataout<=36'h624fd47df;
			11'h6e0: dataout<=36'h1b225f45b;
			11'h6e1: dataout<=36'h3508dd1f8;
			11'h6e2: dataout<=36'h4c8619a67;
			11'h6e3: dataout<=36'h608a15031;
			11'h6e4: dataout<=36'h1a775f4ee;
			11'h6e5: dataout<=36'h33c9dd436;
			11'h6e6: dataout<=36'h4adf19f41;
			11'h6e7: dataout<=36'h5eb8d585d;
			11'h6e8: dataout<=36'h19cbdf57d;
			11'h6e9: dataout<=36'h32889d666;
			11'h6ea: dataout<=36'h49325a401;
			11'h6eb: dataout<=36'h5cdc96060;
			11'h6ec: dataout<=36'h19209f608;
			11'h6ed: dataout<=36'h3146dd887;
			11'h6ee: dataout<=36'h47821a8a2;
			11'h6ef: dataout<=36'h5af59683a;
			11'h6f0: dataout<=36'h1874df690;
			11'h6f1: dataout<=36'h3002dda9c;
			11'h6f2: dataout<=36'h45cc1ad2b;
			11'h6f3: dataout<=36'h590416fea;
			11'h6f4: dataout<=36'h17c91f713;
			11'h6f5: dataout<=36'h2ebdddca0;
			11'h6f6: dataout<=36'h4411db193;
			11'h6f7: dataout<=36'h57081776f;
			11'h6f8: dataout<=36'h171d1f794;
			11'h6f9: dataout<=36'h2d779de9a;
			11'h6fa: dataout<=36'h42535b5e4;
			11'h6fb: dataout<=36'h5501d7ec9;
			11'h6fc: dataout<=36'h1670df810;
			11'h6fd: dataout<=36'h2c2f9e083;
			11'h6fe: dataout<=36'h408fdba14;
			11'h6ff: dataout<=36'h52f1985f5;
			11'h700: dataout<=36'h15c49f889;
			11'h701: dataout<=36'h2ae6de260;
			11'h702: dataout<=36'h3ec91be29;
			11'h703: dataout<=36'h50d7d8cf4;
			11'h704: dataout<=36'h15181f8fe;
			11'h705: dataout<=36'h299c5e42d;
			11'h706: dataout<=36'h3cfd5c21f;
			11'h707: dataout<=36'h4eb4993c5;
			11'h708: dataout<=36'h146b5f970;
			11'h709: dataout<=36'h2850de5ee;
			11'h70a: dataout<=36'h3b2ddc5fa;
			11'h70b: dataout<=36'h4c8819a66;
			11'h70c: dataout<=36'h13be9f9de;
			11'h70d: dataout<=36'h27041e7a0;
			11'h70e: dataout<=36'h395a9c9b6;
			11'h70f: dataout<=36'h4a52da0d8;
			11'h710: dataout<=36'h13119fa48;
			11'h711: dataout<=36'h25b61e944;
			11'h712: dataout<=36'h37831cd54;
			11'h713: dataout<=36'h48149a719;
			11'h714: dataout<=36'h12649faae;
			11'h715: dataout<=36'h24675ead8;
			11'h716: dataout<=36'h35a89d0d2;
			11'h717: dataout<=36'h45ce5ad29;
			11'h718: dataout<=36'h11b75fb11;
			11'h719: dataout<=36'h23175ec60;
			11'h71a: dataout<=36'h33ca5d434;
			11'h71b: dataout<=36'h437f9b306;
			11'h71c: dataout<=36'h110a1fb70;
			11'h71d: dataout<=36'h21c69edd8;
			11'h71e: dataout<=36'h31e91d776;
			11'h71f: dataout<=36'h41291b8b1;
			11'h720: dataout<=36'h105c9fbcb;
			11'h721: dataout<=36'h20745ef42;
			11'h722: dataout<=36'h3003dda98;
			11'h723: dataout<=36'h3ecb1be28;
			11'h724: dataout<=36'h0faf1fc23;
			11'h725: dataout<=36'h1f219f09e;
			11'h726: dataout<=36'h2e1c1dd9d;
			11'h727: dataout<=36'h3c659c36b;
			11'h728: dataout<=36'h0f015fc77;
			11'h729: dataout<=36'h1dcd9f1eb;
			11'h72a: dataout<=36'h2c309e082;
			11'h72b: dataout<=36'h39f91c879;
			11'h72c: dataout<=36'h0e539fcc7;
			11'h72d: dataout<=36'h1c791f32a;
			11'h72e: dataout<=36'h2a42de347;
			11'h72f: dataout<=36'h3785dcd52;
			11'h730: dataout<=36'h0da59fd13;
			11'h731: dataout<=36'h1b235f459;
			11'h732: dataout<=36'h2851de5eb;
			11'h733: dataout<=36'h350c1d1f6;
			11'h734: dataout<=36'h0cf79fd5c;
			11'h735: dataout<=36'h19cd1f57b;
			11'h736: dataout<=36'h265e9e871;
			11'h737: dataout<=36'h328c1d662;
			11'h738: dataout<=36'h0c499fda1;
			11'h739: dataout<=36'h18761f68d;
			11'h73a: dataout<=36'h24689ead5;
			11'h73b: dataout<=36'h30065da98;
			11'h73c: dataout<=36'h0b9b5fde2;
			11'h73d: dataout<=36'h171e1f791;
			11'h73e: dataout<=36'h22701ed1a;
			11'h73f: dataout<=36'h2d7adde97;
			11'h740: dataout<=36'h0aed1fe20;
			11'h741: dataout<=36'h15c5df887;
			11'h742: dataout<=36'h2075def3f;
			11'h743: dataout<=36'h2aea1e25d;
			11'h744: dataout<=36'h0a3e9fe5a;
			11'h745: dataout<=36'h146c5f96e;
			11'h746: dataout<=36'h1e789f144;
			11'h747: dataout<=36'h28545e5ec;
			11'h748: dataout<=36'h09905fe90;
			11'h749: dataout<=36'h13131fa46;
			11'h74a: dataout<=36'h1c7a5f327;
			11'h74b: dataout<=36'h25b9de941;
			11'h74c: dataout<=36'h08e1dfec2;
			11'h74d: dataout<=36'h11b89fb0e;
			11'h74e: dataout<=36'h1a799f4e8;
			11'h74f: dataout<=36'h231adec5e;
			11'h750: dataout<=36'h08331fef1;
			11'h751: dataout<=36'h105d9fbc9;
			11'h752: dataout<=36'h1876df68b;
			11'h753: dataout<=36'h2077def41;
			11'h754: dataout<=36'h07849ff1c;
			11'h755: dataout<=36'h0f029fc75;
			11'h756: dataout<=36'h16735f80c;
			11'h757: dataout<=36'h1dd11f1ea;
			11'h758: dataout<=36'h06d5dff43;
			11'h759: dataout<=36'h0da69fd11;
			11'h75a: dataout<=36'h146d5f96b;
			11'h75b: dataout<=36'h1b26df459;
			11'h75c: dataout<=36'h06271ff67;
			11'h75d: dataout<=36'h0c4a9fda0;
			11'h75e: dataout<=36'h1266dfaab;
			11'h75f: dataout<=36'h18795f68d;
			11'h760: dataout<=36'h05785ff87;
			11'h761: dataout<=36'h0aee1fe1f;
			11'h762: dataout<=36'h105edfbc9;
			11'h763: dataout<=36'h15c91f887;
			11'h764: dataout<=36'h04c99ffa3;
			11'h765: dataout<=36'h09919fe8f;
			11'h766: dataout<=36'h0e561fcc4;
			11'h767: dataout<=36'h13165fa46;
			11'h768: dataout<=36'h041adffbb;
			11'h769: dataout<=36'h08349fef0;
			11'h76a: dataout<=36'h0c4c1fd9e;
			11'h76b: dataout<=36'h10615fbca;
			11'h76c: dataout<=36'h036bdffd0;
			11'h76d: dataout<=36'h06d71ff43;
			11'h76e: dataout<=36'h0a411fe58;
			11'h76f: dataout<=36'h0daa5fd12;
			11'h770: dataout<=36'h02bcdffe0;
			11'h771: dataout<=36'h05795ff85;
			11'h772: dataout<=36'h08355feee;
			11'h773: dataout<=36'h0af19fe20;
			11'h774: dataout<=36'h020e1ffee;
			11'h775: dataout<=36'h041c1ffbb;
			11'h776: dataout<=36'h0629dff66;
			11'h777: dataout<=36'h0837dfef1;
			11'h778: dataout<=36'h015f1fff7;
			11'h779: dataout<=36'h02be1ffdf;
			11'h77a: dataout<=36'h041d1ffb8;
			11'h77b: dataout<=36'h057d1ff87;
			11'h77c: dataout<=36'h015f1fff7;
			11'h77d: dataout<=36'h02be1ffdf;
			11'h77e: dataout<=36'h041d1ffb8;
			11'h77f: dataout<=36'h057d1ff87;
			11'h780: dataout<=36'h000000000;
			11'h781: dataout<=36'h000000000;
			11'h782: dataout<=36'h000000000;
			11'h783: dataout<=36'h000000000;
			11'h784: dataout<=36'h000000000;
			11'h785: dataout<=36'h000000000;
			11'h786: dataout<=36'h000000000;
			11'h787: dataout<=36'h000000000;
			11'h788: dataout<=36'h000000000;
			11'h789: dataout<=36'h000000000;
			11'h78a: dataout<=36'h000000000;
			11'h78b: dataout<=36'h000000000;
			11'h78c: dataout<=36'h000000000;
			11'h78d: dataout<=36'h000000000;
			11'h78e: dataout<=36'h000000000;
			11'h78f: dataout<=36'h000000000;
			11'h790: dataout<=36'h000000000;
			11'h791: dataout<=36'h000000000;
			11'h792: dataout<=36'h000000000;
			11'h793: dataout<=36'h000000000;
			11'h794: dataout<=36'h000000000;
			11'h795: dataout<=36'h000000000;
			11'h796: dataout<=36'h000000000;
			11'h797: dataout<=36'h000000000;
			11'h798: dataout<=36'h000000000;
			11'h799: dataout<=36'h000000000;
			11'h79a: dataout<=36'h000000000;
			11'h79b: dataout<=36'h000000000;
			11'h79c: dataout<=36'h000000000;
			11'h79d: dataout<=36'h000000000;
			11'h79e: dataout<=36'h000000000;
			11'h79f: dataout<=36'h000000000;
			11'h7a0: dataout<=36'h000000000;
			11'h7a1: dataout<=36'h000000000;
			11'h7a2: dataout<=36'h000000000;
			11'h7a3: dataout<=36'h000000000;
			11'h7a4: dataout<=36'h000000000;
			11'h7a5: dataout<=36'h000000000;
			11'h7a6: dataout<=36'h000000000;
			11'h7a7: dataout<=36'h000000000;
			11'h7a8: dataout<=36'h000000000;
			11'h7a9: dataout<=36'h000000000;
			11'h7aa: dataout<=36'h000000000;
			11'h7ab: dataout<=36'h000000000;
			11'h7ac: dataout<=36'h000000000;
			11'h7ad: dataout<=36'h000000000;
			11'h7ae: dataout<=36'h000000000;
			11'h7af: dataout<=36'h000000000;
			11'h7b0: dataout<=36'h000000000;
			11'h7b1: dataout<=36'h000000000;
			11'h7b2: dataout<=36'h000000000;
			11'h7b3: dataout<=36'h000000000;
			11'h7b4: dataout<=36'h000000000;
			11'h7b5: dataout<=36'h000000000;
			11'h7b6: dataout<=36'h000000000;
			11'h7b7: dataout<=36'h000000000;
			11'h7b8: dataout<=36'h000000000;
			11'h7b9: dataout<=36'h000000000;
			11'h7ba: dataout<=36'h000000000;
			11'h7bb: dataout<=36'h000000000;
			11'h7bc: dataout<=36'h000000000;
			11'h7bd: dataout<=36'h000000000;
			11'h7be: dataout<=36'h000000000;
			11'h7bf: dataout<=36'h000000000;
			11'h7c0: dataout<=36'h000000000;
			11'h7c1: dataout<=36'h000000000;
			11'h7c2: dataout<=36'h000000000;
			11'h7c3: dataout<=36'h000000000;
			11'h7c4: dataout<=36'h000000000;
			11'h7c5: dataout<=36'h000000000;
			11'h7c6: dataout<=36'h000000000;
			11'h7c7: dataout<=36'h000000000;
			11'h7c8: dataout<=36'h000000000;
			11'h7c9: dataout<=36'h000000000;
			11'h7ca: dataout<=36'h000000000;
			11'h7cb: dataout<=36'h000000000;
			11'h7cc: dataout<=36'h000000000;
			11'h7cd: dataout<=36'h000000000;
			11'h7ce: dataout<=36'h000000000;
			11'h7cf: dataout<=36'h000000000;
			11'h7d0: dataout<=36'h000000000;
			11'h7d1: dataout<=36'h000000000;
			11'h7d2: dataout<=36'h000000000;
			11'h7d3: dataout<=36'h000000000;
			11'h7d4: dataout<=36'h000000000;
			11'h7d5: dataout<=36'h000000000;
			11'h7d6: dataout<=36'h000000000;
			11'h7d7: dataout<=36'h000000000;
			11'h7d8: dataout<=36'h000000000;
			11'h7d9: dataout<=36'h000000000;
			11'h7da: dataout<=36'h000000000;
			11'h7db: dataout<=36'h000000000;
			11'h7dc: dataout<=36'h000000000;
			11'h7dd: dataout<=36'h000000000;
			11'h7de: dataout<=36'h000000000;
			11'h7df: dataout<=36'h000000000;
			11'h7e0: dataout<=36'h000000000;
			11'h7e1: dataout<=36'h000000000;
			11'h7e2: dataout<=36'h000000000;
			11'h7e3: dataout<=36'h000000000;
			11'h7e4: dataout<=36'h000000000;
			11'h7e5: dataout<=36'h000000000;
			11'h7e6: dataout<=36'h000000000;
			11'h7e7: dataout<=36'h000000000;
			11'h7e8: dataout<=36'h000000000;
			11'h7e9: dataout<=36'h000000000;
			11'h7ea: dataout<=36'h000000000;
			11'h7eb: dataout<=36'h000000000;
			11'h7ec: dataout<=36'h000000000;
			11'h7ed: dataout<=36'h000000000;
			11'h7ee: dataout<=36'h000000000;
			11'h7ef: dataout<=36'h000000000;
			11'h7f0: dataout<=36'h000000000;
			11'h7f1: dataout<=36'h000000000;
			11'h7f2: dataout<=36'h000000000;
			11'h7f3: dataout<=36'h000000000;
			11'h7f4: dataout<=36'h000000000;
			11'h7f5: dataout<=36'h000000000;
			11'h7f6: dataout<=36'h000000000;
			11'h7f7: dataout<=36'h000000000;
			11'h7f8: dataout<=36'h000000000;
			11'h7f9: dataout<=36'h000000000;
			11'h7fa: dataout<=36'h000000000;
			11'h7fb: dataout<=36'h000000000;
			11'h7fc: dataout<=36'h000000000;
			11'h7fd: dataout<=36'h000000000;
			11'h7fe: dataout<=36'h000000000;
			11'h7ff: dataout<=36'h000000000;
		endcase
	end
endmodule

