module nco_rom_4ch_fc2400_fs11718 (clock,addr,dataout);
	input clock;
	input [10:0] addr;
	output reg signed [35:0] dataout;
	always @(posedge clock) begin
		case (addr)
			11'h000: dataout<=36'h7aad49217;
			11'h001: dataout<=36'h460225361;
			11'h002: dataout<=36'had46a794f;
			11'h003: dataout<=36'h8ac7ccda8;
			11'h004: dataout<=36'h7a9449366;
			11'h005: dataout<=36'h4694654e1;
			11'h006: dataout<=36'hae0f676ab;
			11'h007: dataout<=36'h8a3d0c8a4;
			11'h008: dataout<=36'h7a7b094b5;
			11'h009: dataout<=36'h472625664;
			11'h00a: dataout<=36'haed9a740e;
			11'h00b: dataout<=36'h89b58c399;
			11'h00c: dataout<=36'h7a6189604;
			11'h00d: dataout<=36'h47b7657eb;
			11'h00e: dataout<=36'hafa567177;
			11'h00f: dataout<=36'h8931cbe89;
			11'h010: dataout<=36'h7a47c9752;
			11'h011: dataout<=36'h4847e5974;
			11'h012: dataout<=36'hb07226ee9;
			11'h013: dataout<=36'h88b14b973;
			11'h014: dataout<=36'h7a2dc98a0;
			11'h015: dataout<=36'h48d7e5b01;
			11'h016: dataout<=36'hb14066c60;
			11'h017: dataout<=36'h88344b458;
			11'h018: dataout<=36'h7a13899ee;
			11'h019: dataout<=36'h496765c91;
			11'h01a: dataout<=36'hb20fe69de;
			11'h01b: dataout<=36'h87bacaf37;
			11'h01c: dataout<=36'h79f949b3c;
			11'h01d: dataout<=36'h49f6e5e23;
			11'h01e: dataout<=36'hb2e0a6760;
			11'h01f: dataout<=36'h8744caa11;
			11'h020: dataout<=36'h79de89c89;
			11'h021: dataout<=36'h4a8525fba;
			11'h022: dataout<=36'hb3b2e64ec;
			11'h023: dataout<=36'h86d24a4e7;
			11'h024: dataout<=36'h79c3c9dd6;
			11'h025: dataout<=36'h4b1326152;
			11'h026: dataout<=36'hb485e627d;
			11'h027: dataout<=36'h866349fb7;
			11'h028: dataout<=36'h79a889f23;
			11'h029: dataout<=36'h4ba0a62ef;
			11'h02a: dataout<=36'hb55b26016;
			11'h02b: dataout<=36'h85f809a83;
			11'h02c: dataout<=36'h798d4a06f;
			11'h02d: dataout<=36'h4c2d6648e;
			11'h02e: dataout<=36'hb630a5db6;
			11'h02f: dataout<=36'h85900954b;
			11'h030: dataout<=36'h7971ca1bb;
			11'h031: dataout<=36'h4cb9a662f;
			11'h032: dataout<=36'hb70765b5c;
			11'h033: dataout<=36'h852bc900e;
			11'h034: dataout<=36'h79560a307;
			11'h035: dataout<=36'h4d45667d5;
			11'h036: dataout<=36'hb7dfe5909;
			11'h037: dataout<=36'h84cb48acc;
			11'h038: dataout<=36'h793a0a453;
			11'h039: dataout<=36'h4dd0e697d;
			11'h03a: dataout<=36'hb8b9656bc;
			11'h03b: dataout<=36'h846e48587;
			11'h03c: dataout<=36'h791dca59e;
			11'h03d: dataout<=36'h4e5b26b28;
			11'h03e: dataout<=36'hb993e5479;
			11'h03f: dataout<=36'h8414c803e;
			11'h040: dataout<=36'h79018a6e9;
			11'h041: dataout<=36'h4ee566cd5;
			11'h042: dataout<=36'hba6f65239;
			11'h043: dataout<=36'h83bec7af1;
			11'h044: dataout<=36'h78e4ca833;
			11'h045: dataout<=36'h4f6ea6e86;
			11'h046: dataout<=36'hbb4c25004;
			11'h047: dataout<=36'h836cc75a1;
			11'h048: dataout<=36'h78c80a97e;
			11'h049: dataout<=36'h4ff7e703a;
			11'h04a: dataout<=36'hbc2a64dd2;
			11'h04b: dataout<=36'h831e0704d;
			11'h04c: dataout<=36'h78ab0aac8;
			11'h04d: dataout<=36'h5080271f0;
			11'h04e: dataout<=36'hbd0924ba9;
			11'h04f: dataout<=36'h82d346af6;
			11'h050: dataout<=36'h788d8ac11;
			11'h051: dataout<=36'h5107673ab;
			11'h052: dataout<=36'hbde9a498b;
			11'h053: dataout<=36'h828c0659b;
			11'h054: dataout<=36'h78700ad5b;
			11'h055: dataout<=36'h518ee7567;
			11'h056: dataout<=36'hbecb2476e;
			11'h057: dataout<=36'h82484603e;
			11'h058: dataout<=36'h78524aea4;
			11'h059: dataout<=36'h521567727;
			11'h05a: dataout<=36'hbfada455c;
			11'h05b: dataout<=36'h820845ade;
			11'h05c: dataout<=36'h78348afed;
			11'h05d: dataout<=36'h529b678e8;
			11'h05e: dataout<=36'hc090a434f;
			11'h05f: dataout<=36'h81cc0557b;
			11'h060: dataout<=36'h78164b135;
			11'h061: dataout<=36'h5320a7aad;
			11'h062: dataout<=36'hc174e414b;
			11'h063: dataout<=36'h819385016;
			11'h064: dataout<=36'h77f7cb27d;
			11'h065: dataout<=36'h53a527c76;
			11'h066: dataout<=36'hc25aa3f4f;
			11'h067: dataout<=36'h815e84aaf;
			11'h068: dataout<=36'h77d94b3c5;
			11'h069: dataout<=36'h542967e40;
			11'h06a: dataout<=36'hc340e3d58;
			11'h06b: dataout<=36'h812d84545;
			11'h06c: dataout<=36'h77ba8b50d;
			11'h06d: dataout<=36'h54ad6800d;
			11'h06e: dataout<=36'hc428a3b67;
			11'h06f: dataout<=36'h810003fd9;
			11'h070: dataout<=36'h779b8b654;
			11'h071: dataout<=36'h5530281dd;
			11'h072: dataout<=36'hc510e3980;
			11'h073: dataout<=36'h80d643a6b;
			11'h074: dataout<=36'h777c0b79a;
			11'h075: dataout<=36'h55b1e83b2;
			11'h076: dataout<=36'hc5faa37a5;
			11'h077: dataout<=36'h80b0034fc;
			11'h078: dataout<=36'h775ccb8e1;
			11'h079: dataout<=36'h5633e8586;
			11'h07a: dataout<=36'hc6e4a35ca;
			11'h07b: dataout<=36'h808dc2f8b;
			11'h07c: dataout<=36'h773d0ba27;
			11'h07d: dataout<=36'h56b4e875f;
			11'h07e: dataout<=36'hc7cfe33f9;
			11'h07f: dataout<=36'h806f02a19;
			11'h080: dataout<=36'h771d0bb6d;
			11'h081: dataout<=36'h57352893b;
			11'h082: dataout<=36'hc8bc63231;
			11'h083: dataout<=36'h8054424a5;
			11'h084: dataout<=36'h76fd0bcb2;
			11'h085: dataout<=36'h57b4e8b18;
			11'h086: dataout<=36'hc9a92306f;
			11'h087: dataout<=36'h803d01f31;
			11'h088: dataout<=36'h76dc8bdf7;
			11'h089: dataout<=36'h5833e8cfa;
			11'h08a: dataout<=36'hca9762eb7;
			11'h08b: dataout<=36'h8029819bb;
			11'h08c: dataout<=36'h76bc0bf3c;
			11'h08d: dataout<=36'h58b268edd;
			11'h08e: dataout<=36'hcb8662d04;
			11'h08f: dataout<=36'h8019c1445;
			11'h090: dataout<=36'h769b4c081;
			11'h091: dataout<=36'h5930a90c4;
			11'h092: dataout<=36'hcc7662b58;
			11'h093: dataout<=36'h800dc0ece;
			11'h094: dataout<=36'h767a4c1c5;
			11'h095: dataout<=36'h59ada92ad;
			11'h096: dataout<=36'hcd67229b5;
			11'h097: dataout<=36'h800580957;
			11'h098: dataout<=36'h76590c308;
			11'h099: dataout<=36'h5a29e9498;
			11'h09a: dataout<=36'hce582281c;
			11'h09b: dataout<=36'h8001003e0;
			11'h09c: dataout<=36'h76378c44c;
			11'h09d: dataout<=36'h5aa5e9688;
			11'h09e: dataout<=36'hcf4b22688;
			11'h09f: dataout<=36'h80007fe69;
			11'h0a0: dataout<=36'h76160c58f;
			11'h0a1: dataout<=36'h5b2129877;
			11'h0a2: dataout<=36'hd03da24fb;
			11'h0a3: dataout<=36'h80037f8f1;
			11'h0a4: dataout<=36'h75f40c6d1;
			11'h0a5: dataout<=36'h5b9b69a6b;
			11'h0a6: dataout<=36'hd13162379;
			11'h0a7: dataout<=36'h800a3f37a;
			11'h0a8: dataout<=36'h75d20c814;
			11'h0a9: dataout<=36'h5c15a9c62;
			11'h0aa: dataout<=36'hd226a21fc;
			11'h0ab: dataout<=36'h80147ee03;
			11'h0ac: dataout<=36'h75afcc955;
			11'h0ad: dataout<=36'h5c8e69e59;
			11'h0ae: dataout<=36'hd31b22089;
			11'h0af: dataout<=36'h8022be88d;
			11'h0b0: dataout<=36'h758d4ca97;
			11'h0b1: dataout<=36'h5d072a055;
			11'h0b2: dataout<=36'hd411a1f1c;
			11'h0b3: dataout<=36'h8034be317;
			11'h0b4: dataout<=36'h756a8cbd8;
			11'h0b5: dataout<=36'h5d7eea253;
			11'h0b6: dataout<=36'hd50861db8;
			11'h0b7: dataout<=36'h804a3dda2;
			11'h0b8: dataout<=36'h75478cd19;
			11'h0b9: dataout<=36'h5df62a454;
			11'h0ba: dataout<=36'hd60021c5b;
			11'h0bb: dataout<=36'h8063bd82e;
			11'h0bc: dataout<=36'h75244ce59;
			11'h0bd: dataout<=36'h5e6c2a657;
			11'h0be: dataout<=36'hd6f861b09;
			11'h0bf: dataout<=36'h8080bd2bb;
			11'h0c0: dataout<=36'h75010cf99;
			11'h0c1: dataout<=36'h5ee22a85c;
			11'h0c2: dataout<=36'hd7f1219bb;
			11'h0c3: dataout<=36'h80a17cd4a;
			11'h0c4: dataout<=36'h74dd8d0d9;
			11'h0c5: dataout<=36'h5f576aa64;
			11'h0c6: dataout<=36'hd8eaa1876;
			11'h0c7: dataout<=36'h80c5fc7da;
			11'h0c8: dataout<=36'h74b9cd218;
			11'h0c9: dataout<=36'h5fcbaac6e;
			11'h0ca: dataout<=36'hd9e4a173a;
			11'h0cb: dataout<=36'h80ee3c26b;
			11'h0cc: dataout<=36'h7495cd357;
			11'h0cd: dataout<=36'h603f6ae7b;
			11'h0ce: dataout<=36'hdadfa1605;
			11'h0cf: dataout<=36'h811a3bcff;
			11'h0d0: dataout<=36'h74718d496;
			11'h0d1: dataout<=36'h60b2ab08b;
			11'h0d2: dataout<=36'hdbdb614d7;
			11'h0d3: dataout<=36'h8149bb794;
			11'h0d4: dataout<=36'h744d0d5d4;
			11'h0d5: dataout<=36'h6124ab29d;
			11'h0d6: dataout<=36'hdcd7613b4;
			11'h0d7: dataout<=36'h817d3b22c;
			11'h0d8: dataout<=36'h74284d712;
			11'h0d9: dataout<=36'h61966b4b3;
			11'h0da: dataout<=36'hddd4a1298;
			11'h0db: dataout<=36'h81b43acc5;
			11'h0dc: dataout<=36'h74038d84f;
			11'h0dd: dataout<=36'h62072b6c8;
			11'h0de: dataout<=36'hded121184;
			11'h0df: dataout<=36'h81eefa762;
			11'h0e0: dataout<=36'h73de8d98c;
			11'h0e1: dataout<=36'h62776b8e1;
			11'h0e2: dataout<=36'hdfcee1077;
			11'h0e3: dataout<=36'h822d3a200;
			11'h0e4: dataout<=36'h73b94dac9;
			11'h0e5: dataout<=36'h62e6ebafd;
			11'h0e6: dataout<=36'he0cd60f72;
			11'h0e7: dataout<=36'h826f79ca2;
			11'h0e8: dataout<=36'h7393cdc05;
			11'h0e9: dataout<=36'h6355abd1b;
			11'h0ea: dataout<=36'he1cc20e77;
			11'h0eb: dataout<=36'h82b539746;
			11'h0ec: dataout<=36'h736e0dd40;
			11'h0ed: dataout<=36'h63c32bf3b;
			11'h0ee: dataout<=36'he2cb20d85;
			11'h0ef: dataout<=36'h82fe791ee;
			11'h0f0: dataout<=36'h73480de7c;
			11'h0f1: dataout<=36'h6430ac15f;
			11'h0f2: dataout<=36'he3cb60c99;
			11'h0f3: dataout<=36'h834bb8c99;
			11'h0f4: dataout<=36'h73220dfb7;
			11'h0f5: dataout<=36'h649d6c383;
			11'h0f6: dataout<=36'he4cb60bb5;
			11'h0f7: dataout<=36'h839c38747;
			11'h0f8: dataout<=36'h72fb8e0f1;
			11'h0f9: dataout<=36'h6508ac5ab;
			11'h0fa: dataout<=36'he5cbe0add;
			11'h0fb: dataout<=36'h83f0b81f8;
			11'h0fc: dataout<=36'h72d50e22b;
			11'h0fd: dataout<=36'h6573ac7d4;
			11'h0fe: dataout<=36'he6cce0a0a;
			11'h0ff: dataout<=36'h844877cae;
			11'h100: dataout<=36'h72ae4e365;
			11'h101: dataout<=36'h65de2ca00;
			11'h102: dataout<=36'he7cea093e;
			11'h103: dataout<=36'h84a437767;
			11'h104: dataout<=36'h72874e49e;
			11'h105: dataout<=36'h66476cc2e;
			11'h106: dataout<=36'he8d06087d;
			11'h107: dataout<=36'h850337224;
			11'h108: dataout<=36'h72604e5d7;
			11'h109: dataout<=36'h66b06ce5d;
			11'h10a: dataout<=36'he9d2607c2;
			11'h10b: dataout<=36'h8565f6ce5;
			11'h10c: dataout<=36'h7238ce710;
			11'h10d: dataout<=36'h6718ad091;
			11'h10e: dataout<=36'head560710;
			11'h10f: dataout<=36'h85cc367ab;
			11'h110: dataout<=36'h72114e848;
			11'h111: dataout<=36'h67802d2c5;
			11'h112: dataout<=36'hebd860665;
			11'h113: dataout<=36'h863636275;
			11'h114: dataout<=36'h71e98e97f;
			11'h115: dataout<=36'h67e66d4fc;
			11'h116: dataout<=36'hecdb605c5;
			11'h117: dataout<=36'h86a3b5d43;
			11'h118: dataout<=36'h71c18eab7;
			11'h119: dataout<=36'h684cad735;
			11'h11a: dataout<=36'heddf6052a;
			11'h11b: dataout<=36'h8714b5816;
			11'h11c: dataout<=36'h71994ebed;
			11'h11d: dataout<=36'h68b12d970;
			11'h11e: dataout<=36'heee2e049c;
			11'h11f: dataout<=36'h8789352ef;
			11'h120: dataout<=36'h7170ced24;
			11'h121: dataout<=36'h6915adbaf;
			11'h122: dataout<=36'hefe7a0414;
			11'h123: dataout<=36'h880134dcc;
			11'h124: dataout<=36'h71484ee5a;
			11'h125: dataout<=36'h69796ddee;
			11'h126: dataout<=36'hf0ec20392;
			11'h127: dataout<=36'h887cb48ae;
			11'h128: dataout<=36'h711f8ef8f;
			11'h129: dataout<=36'h69dbee02f;
			11'h12a: dataout<=36'hf1f06031b;
			11'h12b: dataout<=36'h88fbb4396;
			11'h12c: dataout<=36'h70f64f0c4;
			11'h12d: dataout<=36'h6a3dae274;
			11'h12e: dataout<=36'hf2f5a02ae;
			11'h12f: dataout<=36'h897e33e84;
			11'h130: dataout<=36'h70cd0f1f9;
			11'h131: dataout<=36'h6a9f2e4ba;
			11'h132: dataout<=36'hf3fb20246;
			11'h133: dataout<=36'h8a0433977;
			11'h134: dataout<=36'h70a3cf32d;
			11'h135: dataout<=36'h6affae701;
			11'h136: dataout<=36'hf500201e7;
			11'h137: dataout<=36'h8a8db346f;
			11'h138: dataout<=36'h707a0f460;
			11'h139: dataout<=36'h6b5eee94b;
			11'h13a: dataout<=36'hf60560193;
			11'h13b: dataout<=36'h8b1a72f6e;
			11'h13c: dataout<=36'h70504f594;
			11'h13d: dataout<=36'h6bbe2eb97;
			11'h13e: dataout<=36'hf70b60143;
			11'h13f: dataout<=36'h8baab2a73;
			11'h140: dataout<=36'h70260f6c7;
			11'h141: dataout<=36'h6c1c2ede6;
			11'h142: dataout<=36'hf811a00ff;
			11'h143: dataout<=36'h8c3e7257e;
			11'h144: dataout<=36'h6ffbcf7f9;
			11'h145: dataout<=36'h6c792f036;
			11'h146: dataout<=36'hf917600c3;
			11'h147: dataout<=36'h8cd572090;
			11'h148: dataout<=36'h6fd14f92b;
			11'h149: dataout<=36'h6cd5af288;
			11'h14a: dataout<=36'hfa1d6008e;
			11'h14b: dataout<=36'h8d6fb1ba7;
			11'h14c: dataout<=36'h6fa6cfa5c;
			11'h14d: dataout<=36'h6d316f4db;
			11'h14e: dataout<=36'hfb2320061;
			11'h14f: dataout<=36'h8e0d716c6;
			11'h150: dataout<=36'h6f7bcfb8d;
			11'h151: dataout<=36'h6d8c2f732;
			11'h152: dataout<=36'hfc29a003f;
			11'h153: dataout<=36'h8eae711ec;
			11'h154: dataout<=36'h6f50cfcbe;
			11'h155: dataout<=36'h6de66f989;
			11'h156: dataout<=36'hfd3020022;
			11'h157: dataout<=36'h8f52f0d18;
			11'h158: dataout<=36'h6f258fdee;
			11'h159: dataout<=36'h6e3fafbe3;
			11'h15a: dataout<=36'hfe366000f;
			11'h15b: dataout<=36'h8ffa7084b;
			11'h15c: dataout<=36'h6efa0ff1d;
			11'h15d: dataout<=36'h6e97efe3e;
			11'h15e: dataout<=36'hff3c60006;
			11'h15f: dataout<=36'h90a570386;
			11'h160: dataout<=36'h6ece5004d;
			11'h161: dataout<=36'h6eeff009d;
			11'h162: dataout<=36'h0043a0003;
			11'h163: dataout<=36'h9153afec8;
			11'h164: dataout<=36'h6ea25017b;
			11'h165: dataout<=36'h6f46702fd;
			11'h166: dataout<=36'h0149e000c;
			11'h167: dataout<=36'h9204efa12;
			11'h168: dataout<=36'h6e76502aa;
			11'h169: dataout<=36'h6f9cf055e;
			11'h16a: dataout<=36'h025060018;
			11'h16b: dataout<=36'h92b9af563;
			11'h16c: dataout<=36'h6e4a103d7;
			11'h16d: dataout<=36'h6ff1f07c0;
			11'h16e: dataout<=36'h035660030;
			11'h16f: dataout<=36'h93716f0bc;
			11'h170: dataout<=36'h6e1d90505;
			11'h171: dataout<=36'h7046b0a26;
			11'h172: dataout<=36'h045d2004e;
			11'h173: dataout<=36'h942c6ec1d;
			11'h174: dataout<=36'h6df0d0631;
			11'h175: dataout<=36'h7099f0c8c;
			11'h176: dataout<=36'h0562e0078;
			11'h177: dataout<=36'h94ea6e786;
			11'h178: dataout<=36'h6dc41075e;
			11'h179: dataout<=36'h70ed30ef4;
			11'h17a: dataout<=36'h0669200a5;
			11'h17b: dataout<=36'h95abae2f7;
			11'h17c: dataout<=36'h6d96d0889;
			11'h17d: dataout<=36'h713e7115f;
			11'h17e: dataout<=36'h076ee00e2;
			11'h17f: dataout<=36'h96702de71;
			11'h180: dataout<=36'h6d69909b5;
			11'h181: dataout<=36'h718ff13cb;
			11'h182: dataout<=36'h087520121;
			11'h183: dataout<=36'h97376d9f3;
			11'h184: dataout<=36'h6d3c10ae0;
			11'h185: dataout<=36'h71e071639;
			11'h186: dataout<=36'h097b2016a;
			11'h187: dataout<=36'h9801ed57d;
			11'h188: dataout<=36'h6d0e50c0a;
			11'h189: dataout<=36'h722fb18a9;
			11'h18a: dataout<=36'h0a80a01bd;
			11'h18b: dataout<=36'h98cf6d110;
			11'h18c: dataout<=36'h6ce090d34;
			11'h18d: dataout<=36'h727e71b19;
			11'h18e: dataout<=36'h0b85e0216;
			11'h18f: dataout<=36'h99a02ccac;
			11'h190: dataout<=36'h6cb250e5d;
			11'h191: dataout<=36'h72cbf1d8c;
			11'h192: dataout<=36'h0c8b2027b;
			11'h193: dataout<=36'h9a73ac851;
			11'h194: dataout<=36'h6c8410f86;
			11'h195: dataout<=36'h7318f2001;
			11'h196: dataout<=36'h0d90602e6;
			11'h197: dataout<=36'h9b4a2c400;
			11'h198: dataout<=36'h6c55910af;
			11'h199: dataout<=36'h736532277;
			11'h19a: dataout<=36'h0e9560358;
			11'h19b: dataout<=36'h9c236bfb7;
			11'h19c: dataout<=36'h6c26d11d6;
			11'h19d: dataout<=36'h73b0324ef;
			11'h19e: dataout<=36'h0f99a03d6;
			11'h19f: dataout<=36'h9cffebb78;
			11'h1a0: dataout<=36'h6bf8112fe;
			11'h1a1: dataout<=36'h73faf2768;
			11'h1a2: dataout<=36'h109e20458;
			11'h1a3: dataout<=36'h9ddf2b742;
			11'h1a4: dataout<=36'h6bc8d1425;
			11'h1a5: dataout<=36'h7444729e4;
			11'h1a6: dataout<=36'h11a2a04e6;
			11'h1a7: dataout<=36'h9ec12b316;
			11'h1a8: dataout<=36'h6b999154b;
			11'h1a9: dataout<=36'h748cf2c5f;
			11'h1aa: dataout<=36'h12a5e057b;
			11'h1ab: dataout<=36'h9fa62aef3;
			11'h1ac: dataout<=36'h6b6a11671;
			11'h1ad: dataout<=36'h74d4f2ede;
			11'h1ae: dataout<=36'h13a9a0618;
			11'h1af: dataout<=36'ha08deaadb;
			11'h1b0: dataout<=36'h6b3a91796;
			11'h1b1: dataout<=36'h751bf315c;
			11'h1b2: dataout<=36'h14ac206bc;
			11'h1b3: dataout<=36'ha1786a6cc;
			11'h1b4: dataout<=36'h6b0a918bb;
			11'h1b5: dataout<=36'h7562333de;
			11'h1b6: dataout<=36'h15af6076b;
			11'h1b7: dataout<=36'ha265aa2c7;
			11'h1b8: dataout<=36'h6ada919e0;
			11'h1b9: dataout<=36'h75a7b3661;
			11'h1ba: dataout<=36'h16b220820;
			11'h1bb: dataout<=36'ha355a9ecd;
			11'h1bc: dataout<=36'h6aaa51b04;
			11'h1bd: dataout<=36'h75ec338e5;
			11'h1be: dataout<=36'h17b4208de;
			11'h1bf: dataout<=36'ha44869add;
			11'h1c0: dataout<=36'h6a79d1c27;
			11'h1c1: dataout<=36'h762fb3b6a;
			11'h1c2: dataout<=36'h18b5a09a5;
			11'h1c3: dataout<=36'ha53de96f7;
			11'h1c4: dataout<=36'h6a4951d4a;
			11'h1c5: dataout<=36'h7672b3df0;
			11'h1c6: dataout<=36'h19b6e0a72;
			11'h1c7: dataout<=36'ha635e931c;
			11'h1c8: dataout<=36'h6a1851e6c;
			11'h1c9: dataout<=36'h76b434079;
			11'h1ca: dataout<=36'h1ab7a0b4b;
			11'h1cb: dataout<=36'ha730a8f4b;
			11'h1cc: dataout<=36'h69e751f8e;
			11'h1cd: dataout<=36'h76f574303;
			11'h1ce: dataout<=36'h1bb860c2a;
			11'h1cf: dataout<=36'ha82de8b86;
			11'h1d0: dataout<=36'h69b6120af;
			11'h1d1: dataout<=36'h77357458e;
			11'h1d2: dataout<=36'h1cb820d12;
			11'h1d3: dataout<=36'ha92da87cb;
			11'h1d4: dataout<=36'h6984921d0;
			11'h1d5: dataout<=36'h7774b481b;
			11'h1d6: dataout<=36'h1db7e0e02;
			11'h1d7: dataout<=36'haa302841b;
			11'h1d8: dataout<=36'h6953122f0;
			11'h1d9: dataout<=36'h77b334aa8;
			11'h1da: dataout<=36'h1eb6a0ef9;
			11'h1db: dataout<=36'hab34e8076;
			11'h1dc: dataout<=36'h692152410;
			11'h1dd: dataout<=36'h77f0f4d37;
			11'h1de: dataout<=36'h1fb560ff7;
			11'h1df: dataout<=36'hac3c67cdd;
			11'h1e0: dataout<=36'h68ef5252f;
			11'h1e1: dataout<=36'h782d74fc7;
			11'h1e2: dataout<=36'h20b321100;
			11'h1e3: dataout<=36'had462794e;
			11'h1e4: dataout<=36'h68bd1264d;
			11'h1e5: dataout<=36'h7868f5259;
			11'h1e6: dataout<=36'h21b061212;
			11'h1e7: dataout<=36'hae52675cb;
			11'h1e8: dataout<=36'h688ad276b;
			11'h1e9: dataout<=36'h78a3f54eb;
			11'h1ea: dataout<=36'h22ad21329;
			11'h1eb: dataout<=36'haf60e7254;
			11'h1ec: dataout<=36'h685812889;
			11'h1ed: dataout<=36'h78ddf5781;
			11'h1ee: dataout<=36'h23a9e144b;
			11'h1ef: dataout<=36'hb071e6ee8;
			11'h1f0: dataout<=36'h6825529a6;
			11'h1f1: dataout<=36'h791735a16;
			11'h1f2: dataout<=36'h24a5a1572;
			11'h1f3: dataout<=36'hb18526b88;
			11'h1f4: dataout<=36'h67f252ac2;
			11'h1f5: dataout<=36'h794f35cad;
			11'h1f6: dataout<=36'h25a0a16a4;
			11'h1f7: dataout<=36'hb29aa6834;
			11'h1f8: dataout<=36'h67bf52bde;
			11'h1f9: dataout<=36'h7986b5f44;
			11'h1fa: dataout<=36'h269b217dc;
			11'h1fb: dataout<=36'hb3b2a64ec;
			11'h1fc: dataout<=36'h678c12cfa;
			11'h1fd: dataout<=36'h79bdb61dd;
			11'h1fe: dataout<=36'h27956191a;
			11'h1ff: dataout<=36'hb4cca61af;
			11'h200: dataout<=36'h675852e14;
			11'h201: dataout<=36'h79f2b6478;
			11'h202: dataout<=36'h288e61a66;
			11'h203: dataout<=36'hb5e8e5e7f;
			11'h204: dataout<=36'h6724d2f2f;
			11'h205: dataout<=36'h7a27f6713;
			11'h206: dataout<=36'h298721bb4;
			11'h207: dataout<=36'hb70725b5b;
			11'h208: dataout<=36'h66f0d3048;
			11'h209: dataout<=36'h7a5b369af;
			11'h20a: dataout<=36'h2a7ea1d0e;
			11'h20b: dataout<=36'hb827a5843;
			11'h20c: dataout<=36'h66bcd3161;
			11'h20d: dataout<=36'h7a8e36c4c;
			11'h20e: dataout<=36'h2b75a1e6e;
			11'h20f: dataout<=36'hb94a65538;
			11'h210: dataout<=36'h66889327a;
			11'h211: dataout<=36'h7ac076eeb;
			11'h212: dataout<=36'h2c6c61fd6;
			11'h213: dataout<=36'hba6f25239;
			11'h214: dataout<=36'h665413392;
			11'h215: dataout<=36'h7af17718b;
			11'h216: dataout<=36'h2d6222147;
			11'h217: dataout<=36'hbb95e4f46;
			11'h218: dataout<=36'h661f534a9;
			11'h219: dataout<=36'h7b217742c;
			11'h21a: dataout<=36'h2e57222c0;
			11'h21b: dataout<=36'hbcbea4c61;
			11'h21c: dataout<=36'h65ea935c0;
			11'h21d: dataout<=36'h7b50f76cd;
			11'h21e: dataout<=36'h2f4b6243f;
			11'h21f: dataout<=36'hbde924988;
			11'h220: dataout<=36'h65b5936d7;
			11'h221: dataout<=36'h7b7fb7970;
			11'h222: dataout<=36'h303f225c6;
			11'h223: dataout<=36'hbf15e46bb;
			11'h224: dataout<=36'h6580537ec;
			11'h225: dataout<=36'h7bacb7c13;
			11'h226: dataout<=36'h313122757;
			11'h227: dataout<=36'hc044643fc;
			11'h228: dataout<=36'h654b13902;
			11'h229: dataout<=36'h7bd9f7eb8;
			11'h22a: dataout<=36'h3223a28ec;
			11'h22b: dataout<=36'hc174a414a;
			11'h22c: dataout<=36'h651553a16;
			11'h22d: dataout<=36'h7c053815e;
			11'h22e: dataout<=36'h331462a8d;
			11'h22f: dataout<=36'hc2a6e3ea4;
			11'h230: dataout<=36'h64df93b2a;
			11'h231: dataout<=36'h7c2ff8405;
			11'h232: dataout<=36'h3404a2c35;
			11'h233: dataout<=36'hc3dae3c0c;
			11'h234: dataout<=36'h64a993c3e;
			11'h235: dataout<=36'h7c59f86ad;
			11'h236: dataout<=36'h34f462de3;
			11'h237: dataout<=36'hc510a3981;
			11'h238: dataout<=36'h647393d51;
			11'h239: dataout<=36'h7c8338955;
			11'h23a: dataout<=36'h35e2e2f98;
			11'h23b: dataout<=36'hc64823703;
			11'h23c: dataout<=36'h643d53e63;
			11'h23d: dataout<=36'h7cab38bfd;
			11'h23e: dataout<=36'h36d023155;
			11'h23f: dataout<=36'hc78163493;
			11'h240: dataout<=36'h6406d3f75;
			11'h241: dataout<=36'h7cd278ea8;
			11'h242: dataout<=36'h37bd2331b;
			11'h243: dataout<=36'hc8bc23230;
			11'h244: dataout<=36'h63d014086;
			11'h245: dataout<=36'h7cf8b9153;
			11'h246: dataout<=36'h38a8e34e8;
			11'h247: dataout<=36'hc9f8a2fda;
			11'h248: dataout<=36'h639954196;
			11'h249: dataout<=36'h7d1df93fd;
			11'h24a: dataout<=36'h3993236bc;
			11'h24b: dataout<=36'hcb3662d92;
			11'h24c: dataout<=36'h6362142a6;
			11'h24d: dataout<=36'h7d42396ab;
			11'h24e: dataout<=36'h3a7d2389a;
			11'h24f: dataout<=36'hcc7622b58;
			11'h250: dataout<=36'h632b143b6;
			11'h251: dataout<=36'h7d6639957;
			11'h252: dataout<=36'h3b6663a7a;
			11'h253: dataout<=36'hcdb72292b;
			11'h254: dataout<=36'h62f3944c5;
			11'h255: dataout<=36'h7d88b9c06;
			11'h256: dataout<=36'h3c4e63c66;
			11'h257: dataout<=36'hcef9a270c;
			11'h258: dataout<=36'h62bc145d3;
			11'h259: dataout<=36'h7daa79eb4;
			11'h25a: dataout<=36'h3d3563e58;
			11'h25b: dataout<=36'hd03da24fb;
			11'h25c: dataout<=36'h6284546e0;
			11'h25d: dataout<=36'h7dcafa163;
			11'h25e: dataout<=36'h3e1ae4052;
			11'h25f: dataout<=36'hd182e22f7;
			11'h260: dataout<=36'h624c547ed;
			11'h261: dataout<=36'h7deafa413;
			11'h262: dataout<=36'h3effe4253;
			11'h263: dataout<=36'hd2c9a2102;
			11'h264: dataout<=36'h6214148fa;
			11'h265: dataout<=36'h7e09fa6c6;
			11'h266: dataout<=36'h3fe46445d;
			11'h267: dataout<=36'hd411a1f1b;
			11'h268: dataout<=36'h61dbd4a06;
			11'h269: dataout<=36'h7e27fa977;
			11'h26a: dataout<=36'h40c72466c;
			11'h26b: dataout<=36'hd55ae1d41;
			11'h26c: dataout<=36'h61a354b11;
			11'h26d: dataout<=36'h7e44fac29;
			11'h26e: dataout<=36'h41a8e4884;
			11'h26f: dataout<=36'hd6a561b76;
			11'h270: dataout<=36'h616ad4c1b;
			11'h271: dataout<=36'h7e613aeda;
			11'h272: dataout<=36'h428924aa0;
			11'h273: dataout<=36'hd7f1219b9;
			11'h274: dataout<=36'h6131d4d25;
			11'h275: dataout<=36'h7e7c3b18e;
			11'h276: dataout<=36'h4368e4cc7;
			11'h277: dataout<=36'hd93e2180a;
			11'h278: dataout<=36'h60f8d4e2f;
			11'h279: dataout<=36'h7e96bb443;
			11'h27a: dataout<=36'h4447e4ef4;
			11'h27b: dataout<=36'hda8c21669;
			11'h27c: dataout<=36'h60bfd4f38;
			11'h27d: dataout<=36'h7eb07b6f6;
			11'h27e: dataout<=36'h452525124;
			11'h27f: dataout<=36'hdbdb214d7;
			11'h280: dataout<=36'h608655040;
			11'h281: dataout<=36'h7ec8bb9ac;
			11'h282: dataout<=36'h460165361;
			11'h283: dataout<=36'hdd2b61353;
			11'h284: dataout<=36'h604cd5147;
			11'h285: dataout<=36'h7ee03bc60;
			11'h286: dataout<=36'h46dc255a2;
			11'h287: dataout<=36'hde7ca11dd;
			11'h288: dataout<=36'h60131524e;
			11'h289: dataout<=36'h7ef6bbf16;
			11'h28a: dataout<=36'h47b6257eb;
			11'h28b: dataout<=36'hdfcee1076;
			11'h28c: dataout<=36'h5fd955355;
			11'h28d: dataout<=36'h7f0cfc1cd;
			11'h28e: dataout<=36'h488f65a39;
			11'h28f: dataout<=36'he121e0f1d;
			11'h290: dataout<=36'h5f9f1545a;
			11'h291: dataout<=36'h7f213c484;
			11'h292: dataout<=36'h496665c92;
			11'h293: dataout<=36'he275e0dd3;
			11'h294: dataout<=36'h5f64d5560;
			11'h295: dataout<=36'h7f357c73c;
			11'h296: dataout<=36'h4a3da5eef;
			11'h297: dataout<=36'he3cae0c97;
			11'h298: dataout<=36'h5f2a95664;
			11'h299: dataout<=36'h7f487c9f3;
			11'h29a: dataout<=36'h4b1266152;
			11'h29b: dataout<=36'he520a0b6a;
			11'h29c: dataout<=36'h5eefd5768;
			11'h29d: dataout<=36'h7f5a3ccac;
			11'h29e: dataout<=36'h4be6663bf;
			11'h29f: dataout<=36'he67720a4b;
			11'h2a0: dataout<=36'h5eb51586b;
			11'h2a1: dataout<=36'h7f6b3cf64;
			11'h2a2: dataout<=36'h4cb8e6630;
			11'h2a3: dataout<=36'he7ce6093b;
			11'h2a4: dataout<=36'h5e7a5596e;
			11'h2a5: dataout<=36'h7f7bbd21c;
			11'h2a6: dataout<=36'h4d8aa68a7;
			11'h2a7: dataout<=36'he9262083a;
			11'h2a8: dataout<=36'h5e3f15a70;
			11'h2a9: dataout<=36'h7f8abd4d6;
			11'h2aa: dataout<=36'h4e5aa6b28;
			11'h2ab: dataout<=36'hea7ee0748;
			11'h2ac: dataout<=36'h5e03d5b71;
			11'h2ad: dataout<=36'h7f98fd78f;
			11'h2ae: dataout<=36'h4f2966dad;
			11'h2af: dataout<=36'hebd820664;
			11'h2b0: dataout<=36'h5dc855c72;
			11'h2b1: dataout<=36'h7fa67da4a;
			11'h2b2: dataout<=36'h4ff76703a;
			11'h2b3: dataout<=36'hed31e058f;
			11'h2b4: dataout<=36'h5d8cd5d72;
			11'h2b5: dataout<=36'h7fb2fdd03;
			11'h2b6: dataout<=36'h50c3672cc;
			11'h2b7: dataout<=36'hee8c604c9;
			11'h2b8: dataout<=36'h5d5115e71;
			11'h2b9: dataout<=36'h7fbe7dfbc;
			11'h2ba: dataout<=36'h518e27565;
			11'h2bb: dataout<=36'hefe720411;
			11'h2bc: dataout<=36'h5d1515f70;
			11'h2bd: dataout<=36'h7fc8fe278;
			11'h2be: dataout<=36'h5257e7806;
			11'h2bf: dataout<=36'hf142a0369;
			11'h2c0: dataout<=36'h5cd8d606e;
			11'h2c1: dataout<=36'h7fd27e533;
			11'h2c2: dataout<=36'h532027aad;
			11'h2c3: dataout<=36'hf29e602cf;
			11'h2c4: dataout<=36'h5c9c9616b;
			11'h2c5: dataout<=36'h7fdafe7ed;
			11'h2c6: dataout<=36'h53e6a7d5a;
			11'h2c7: dataout<=36'hf3faa0244;
			11'h2c8: dataout<=36'h5c6016268;
			11'h2c9: dataout<=36'h7fe2beaa8;
			11'h2ca: dataout<=36'h54ac2800d;
			11'h2cb: dataout<=36'hf557201c8;
			11'h2cc: dataout<=36'h5c2396365;
			11'h2cd: dataout<=36'h7fe9fed64;
			11'h2ce: dataout<=36'h5570a82c6;
			11'h2cf: dataout<=36'hf6b3e015b;
			11'h2d0: dataout<=36'h5be696460;
			11'h2d1: dataout<=36'h7fef7f020;
			11'h2d2: dataout<=36'h563328588;
			11'h2d3: dataout<=36'hf811200fd;
			11'h2d4: dataout<=36'h5ba9d655b;
			11'h2d5: dataout<=36'h7ff4bf2da;
			11'h2d6: dataout<=36'h56f46884b;
			11'h2d7: dataout<=36'hf96e600ad;
			11'h2d8: dataout<=36'h5b6c96655;
			11'h2d9: dataout<=36'h7ff87f596;
			11'h2da: dataout<=36'h57b428b19;
			11'h2db: dataout<=36'hfacbe006d;
			11'h2dc: dataout<=36'h5b2f5674f;
			11'h2dd: dataout<=36'h7ffbff852;
			11'h2de: dataout<=36'h5872e8dea;
			11'h2df: dataout<=36'hfc29a003b;
			11'h2e0: dataout<=36'h5af1d6848;
			11'h2e1: dataout<=36'h7ffdffb0e;
			11'h2e2: dataout<=36'h592fe90c3;
			11'h2e3: dataout<=36'hfd8760019;
			11'h2e4: dataout<=36'h5ab416940;
			11'h2e5: dataout<=36'h7ffeffdca;
			11'h2e6: dataout<=36'h59eb293a3;
			11'h2e7: dataout<=36'hfee560005;
			11'h2e8: dataout<=36'h5a7656a38;
			11'h2e9: dataout<=36'h7fff40086;
			11'h2ea: dataout<=36'h5aa569686;
			11'h2eb: dataout<=36'h0042e0001;
			11'h2ec: dataout<=36'h5a3856b2f;
			11'h2ed: dataout<=36'h7ffe80342;
			11'h2ee: dataout<=36'h5b5de9971;
			11'h2ef: dataout<=36'h01a0e000b;
			11'h2f0: dataout<=36'h59fa56c25;
			11'h2f1: dataout<=36'h7ffd005fc;
			11'h2f2: dataout<=36'h5c14a9c60;
			11'h2f3: dataout<=36'h02fea0024;
			11'h2f4: dataout<=36'h59bbd6d1b;
			11'h2f5: dataout<=36'h7ffa808ba;
			11'h2f6: dataout<=36'h5ccaa9f58;
			11'h2f7: dataout<=36'h045c6004d;
			11'h2f8: dataout<=36'h597d96e10;
			11'h2f9: dataout<=36'h7ff740b74;
			11'h2fa: dataout<=36'h5d7e6a251;
			11'h2fb: dataout<=36'h05ba20084;
			11'h2fc: dataout<=36'h593ed6f04;
			11'h2fd: dataout<=36'h7ff280e30;
			11'h2fe: dataout<=36'h5e30aa555;
			11'h2ff: dataout<=36'h0717a00ca;
			11'h300: dataout<=36'h590016ff8;
			11'h301: dataout<=36'h7fed810ec;
			11'h302: dataout<=36'h5ee1ea85b;
			11'h303: dataout<=36'h0874e011f;
			11'h304: dataout<=36'h58c1170eb;
			11'h305: dataout<=36'h7fe7413a8;
			11'h306: dataout<=36'h5f916ab69;
			11'h307: dataout<=36'h09d1e0183;
			11'h308: dataout<=36'h5882171dd;
			11'h309: dataout<=36'h7fe001662;
			11'h30a: dataout<=36'h603eeae7a;
			11'h30b: dataout<=36'h0b2ea01f6;
			11'h30c: dataout<=36'h5842d72ce;
			11'h30d: dataout<=36'h7fd7c191c;
			11'h30e: dataout<=36'h60eaab192;
			11'h30f: dataout<=36'h0c8ae0277;
			11'h310: dataout<=36'h5803573bf;
			11'h311: dataout<=36'h7fce81bd7;
			11'h312: dataout<=36'h61952b4b0;
			11'h313: dataout<=36'h0de720308;
			11'h314: dataout<=36'h57c3974b0;
			11'h315: dataout<=36'h7fc4c1e94;
			11'h316: dataout<=36'h623eeb7d5;
			11'h317: dataout<=36'h0f42a03a7;
			11'h318: dataout<=36'h5783d759f;
			11'h319: dataout<=36'h7fb98214d;
			11'h31a: dataout<=36'h62e5abafd;
			11'h31b: dataout<=36'h109de0456;
			11'h31c: dataout<=36'h57441768e;
			11'h31d: dataout<=36'h7fae02407;
			11'h31e: dataout<=36'h638bebe29;
			11'h31f: dataout<=36'h11f8a0513;
			11'h320: dataout<=36'h5703d777c;
			11'h321: dataout<=36'h7fa0c26c1;
			11'h322: dataout<=36'h642f6c15e;
			11'h323: dataout<=36'h1352a05df;
			11'h324: dataout<=36'h56c3d786a;
			11'h325: dataout<=36'h7f93c297a;
			11'h326: dataout<=36'h64d2ac493;
			11'h327: dataout<=36'h14ac606b9;
			11'h328: dataout<=36'h568357957;
			11'h329: dataout<=36'h7f8502c35;
			11'h32a: dataout<=36'h6573ac7d3;
			11'h32b: dataout<=36'h1605607a3;
			11'h32c: dataout<=36'h5642d7a43;
			11'h32d: dataout<=36'h7f7542eed;
			11'h32e: dataout<=36'h66126cb15;
			11'h32f: dataout<=36'h175da089b;
			11'h330: dataout<=36'h560217b2e;
			11'h331: dataout<=36'h7f64c31a5;
			11'h332: dataout<=36'h66aface5c;
			11'h333: dataout<=36'h18b5609a2;
			11'h334: dataout<=36'h55c117c19;
			11'h335: dataout<=36'h7f530345f;
			11'h336: dataout<=36'h674bad1ab;
			11'h337: dataout<=36'h1a0c60ab7;
			11'h338: dataout<=36'h558017d03;
			11'h339: dataout<=36'h7f40c3717;
			11'h33a: dataout<=36'h67e5ed4fd;
			11'h33b: dataout<=36'h1b62a0bdb;
			11'h33c: dataout<=36'h553f17ded;
			11'h33d: dataout<=36'h7f2e039ce;
			11'h33e: dataout<=36'h687ead851;
			11'h33f: dataout<=36'h1cb7e0d0e;
			11'h340: dataout<=36'h54fd97ed5;
			11'h341: dataout<=36'h7f1943c85;
			11'h342: dataout<=36'h6914edbae;
			11'h343: dataout<=36'h1e0ca0e4f;
			11'h344: dataout<=36'h54bc17fbd;
			11'h345: dataout<=36'h7f0403f3c;
			11'h346: dataout<=36'h69a9adf0f;
			11'h347: dataout<=36'h1f6020f9f;
			11'h348: dataout<=36'h547a980a5;
			11'h349: dataout<=36'h7eee841f2;
			11'h34a: dataout<=36'h6a3dae271;
			11'h34b: dataout<=36'h20b2e10fe;
			11'h34c: dataout<=36'h5438d818b;
			11'h34d: dataout<=36'h7ed7444a7;
			11'h34e: dataout<=36'h6aceae5db;
			11'h34f: dataout<=36'h2204e126a;
			11'h350: dataout<=36'h53f6d8271;
			11'h351: dataout<=36'h7ebf4475d;
			11'h352: dataout<=36'h6b5e6e94a;
			11'h353: dataout<=36'h2355a13e6;
			11'h354: dataout<=36'h53b498356;
			11'h355: dataout<=36'h7ea644a12;
			11'h356: dataout<=36'h6bec2ecbe;
			11'h357: dataout<=36'h24a56156f;
			11'h358: dataout<=36'h53725843b;
			11'h359: dataout<=36'h7e8c84cc7;
			11'h35a: dataout<=36'h6c78af036;
			11'h35b: dataout<=36'h25f421707;
			11'h35c: dataout<=36'h53301851e;
			11'h35d: dataout<=36'h7e7204f78;
			11'h35e: dataout<=36'h6d02af3af;
			11'h35f: dataout<=36'h2741a18ad;
			11'h360: dataout<=36'h52ed98602;
			11'h361: dataout<=36'h7e56c522d;
			11'h362: dataout<=36'h6d8c2f72f;
			11'h363: dataout<=36'h288e21a61;
			11'h364: dataout<=36'h52aad86e4;
			11'h365: dataout<=36'h7e3a054df;
			11'h366: dataout<=36'h6e12afab4;
			11'h367: dataout<=36'h29d961c24;
			11'h368: dataout<=36'h5267d87c5;
			11'h369: dataout<=36'h7e1c05790;
			11'h36a: dataout<=36'h6e972fe3e;
			11'h36b: dataout<=36'h2b23a1df5;
			11'h36c: dataout<=36'h5224d88a6;
			11'h36d: dataout<=36'h7dfdc5a42;
			11'h36e: dataout<=36'h6f1a701cc;
			11'h36f: dataout<=36'h2c6c61fd3;
			11'h370: dataout<=36'h51e1d8987;
			11'h371: dataout<=36'h7ddf05cf2;
			11'h372: dataout<=36'h6f9c7055b;
			11'h373: dataout<=36'h2db3e21c0;
			11'h374: dataout<=36'h519e58a66;
			11'h375: dataout<=36'h7dbe45fa2;
			11'h376: dataout<=36'h701b708f2;
			11'h377: dataout<=36'h2efa223bb;
			11'h378: dataout<=36'h515ad8b45;
			11'h379: dataout<=36'h7d9d46252;
			11'h37a: dataout<=36'h709970c8c;
			11'h37b: dataout<=36'h303ee25c3;
			11'h37c: dataout<=36'h511758c23;
			11'h37d: dataout<=36'h7d7b46500;
			11'h37e: dataout<=36'h711571028;
			11'h37f: dataout<=36'h3182227da;
			11'h380: dataout<=36'h50d398d00;
			11'h381: dataout<=36'h7d58467ad;
			11'h382: dataout<=36'h718f313c9;
			11'h383: dataout<=36'h32c4229fe;
			11'h384: dataout<=36'h508f98ddd;
			11'h385: dataout<=36'h7d3446a5b;
			11'h386: dataout<=36'h720771770;
			11'h387: dataout<=36'h3404a2c30;
			11'h388: dataout<=36'h504b98eb9;
			11'h389: dataout<=36'h7d0fc6d07;
			11'h38a: dataout<=36'h727df1b18;
			11'h38b: dataout<=36'h3543a2e70;
			11'h38c: dataout<=36'h500758f94;
			11'h38d: dataout<=36'h7ce9c6fb3;
			11'h38e: dataout<=36'h72f231ec6;
			11'h38f: dataout<=36'h3680e30bd;
			11'h390: dataout<=36'h4fc31906e;
			11'h391: dataout<=36'h7cc34725c;
			11'h392: dataout<=36'h736472275;
			11'h393: dataout<=36'h37bce3318;
			11'h394: dataout<=36'h4f7e99148;
			11'h395: dataout<=36'h7c9bc7506;
			11'h396: dataout<=36'h73d532629;
			11'h397: dataout<=36'h38f6e3580;
			11'h398: dataout<=36'h4f3a19221;
			11'h399: dataout<=36'h7c73877af;
			11'h39a: dataout<=36'h7444329e0;
			11'h39b: dataout<=36'h3a2f637f6;
			11'h39c: dataout<=36'h4ef5192f9;
			11'h39d: dataout<=36'h7c49c7a57;
			11'h39e: dataout<=36'h74b072d9d;
			11'h39f: dataout<=36'h3b6663a78;
			11'h3a0: dataout<=36'h4eb0593d1;
			11'h3a1: dataout<=36'h7c2007cff;
			11'h3a2: dataout<=36'h751c3315b;
			11'h3a3: dataout<=36'h3c9b63d09;
			11'h3a4: dataout<=36'h4e6b194a7;
			11'h3a5: dataout<=36'h7bf447fa4;
			11'h3a6: dataout<=36'h75843351e;
			11'h3a7: dataout<=36'h3dcea3fa6;
			11'h3a8: dataout<=36'h4e261957d;
			11'h3a9: dataout<=36'h7bc888249;
			11'h3aa: dataout<=36'h75eb738e2;
			11'h3ab: dataout<=36'h3f0024250;
			11'h3ac: dataout<=36'h4de099653;
			11'h3ad: dataout<=36'h7b9b884ef;
			11'h3ae: dataout<=36'h7650f3cad;
			11'h3af: dataout<=36'h402fe4508;
			11'h3b0: dataout<=36'h4d9b19727;
			11'h3b1: dataout<=36'h7b6d88791;
			11'h3b2: dataout<=36'h76b3b4078;
			11'h3b3: dataout<=36'h415da47cc;
			11'h3b4: dataout<=36'h4d55997fb;
			11'h3b5: dataout<=36'h7b3f08a33;
			11'h3b6: dataout<=36'h771534445;
			11'h3b7: dataout<=36'h4289a4a9d;
			11'h3b8: dataout<=36'h4d0fd98ce;
			11'h3b9: dataout<=36'h7b0f48cd5;
			11'h3ba: dataout<=36'h777474818;
			11'h3bb: dataout<=36'h43b364d7b;
			11'h3bc: dataout<=36'h4cc9d99a0;
			11'h3bd: dataout<=36'h7ade88f75;
			11'h3be: dataout<=36'h77d174bee;
			11'h3bf: dataout<=36'h44db65066;
			11'h3c0: dataout<=36'h4c83d9a72;
			11'h3c1: dataout<=36'h7aad49214;
			11'h3c2: dataout<=36'h782cf4fc5;
			11'h3c3: dataout<=36'h46016535d;
			11'h3c4: dataout<=36'h4c3d99b43;
			11'h3c5: dataout<=36'h7a7b094b3;
			11'h3c6: dataout<=36'h7886b53a0;
			11'h3c7: dataout<=36'h472565661;
			11'h3c8: dataout<=36'h4bf759c13;
			11'h3c9: dataout<=36'h7a47c9750;
			11'h3ca: dataout<=36'h78ddf577e;
			11'h3cb: dataout<=36'h484725971;
			11'h3cc: dataout<=36'h4bb0d9ce2;
			11'h3cd: dataout<=36'h7a13899eb;
			11'h3ce: dataout<=36'h7932f5b5e;
			11'h3cf: dataout<=36'h4966e5c8d;
			11'h3d0: dataout<=36'h4b6a19db0;
			11'h3d1: dataout<=36'h79de09c86;
			11'h3d2: dataout<=36'h7985f5f43;
			11'h3d3: dataout<=36'h4a8465fb6;
			11'h3d4: dataout<=36'h4b2359e7e;
			11'h3d5: dataout<=36'h79a849f20;
			11'h3d6: dataout<=36'h79d776329;
			11'h3d7: dataout<=36'h4b9fe62eb;
			11'h3d8: dataout<=36'h4adc99f4b;
			11'h3d9: dataout<=36'h79718a1b8;
			11'h3da: dataout<=36'h7a26f6710;
			11'h3db: dataout<=36'h4cb92662c;
			11'h3dc: dataout<=36'h4a959a017;
			11'h3dd: dataout<=36'h7939ca44f;
			11'h3de: dataout<=36'h7a7436afb;
			11'h3df: dataout<=36'h4dd026979;
			11'h3e0: dataout<=36'h4a4e5a0e3;
			11'h3e1: dataout<=36'h79014a6e6;
			11'h3e2: dataout<=36'h7abfb6ee9;
			11'h3e3: dataout<=36'h4ee4a6cd1;
			11'h3e4: dataout<=36'h4a071a1ae;
			11'h3e5: dataout<=36'h78c80a97c;
			11'h3e6: dataout<=36'h7b09772d9;
			11'h3e7: dataout<=36'h4ff727036;
			11'h3e8: dataout<=36'h49bf9a278;
			11'h3e9: dataout<=36'h788d8ac10;
			11'h3ea: dataout<=36'h7b50b76cc;
			11'h3eb: dataout<=36'h5107273a6;
			11'h3ec: dataout<=36'h49781a341;
			11'h3ed: dataout<=36'h78524aea1;
			11'h3ee: dataout<=36'h7b95f7abf;
			11'h3ef: dataout<=36'h5214e7722;
			11'h3f0: dataout<=36'h49305a409;
			11'h3f1: dataout<=36'h78160b132;
			11'h3f2: dataout<=36'h7bd8f7eb6;
			11'h3f3: dataout<=36'h532027aa9;
			11'h3f4: dataout<=36'h48e89a4d1;
			11'h3f5: dataout<=36'h77d94b3c2;
			11'h3f6: dataout<=36'h7c1a782ae;
			11'h3f7: dataout<=36'h542927e3c;
			11'h3f8: dataout<=36'h48a09a598;
			11'h3f9: dataout<=36'h779b4b651;
			11'h3fa: dataout<=36'h7c59b86a9;
			11'h3fb: dataout<=36'h552f681da;
			11'h3fc: dataout<=36'h48585a65e;
			11'h3fd: dataout<=36'h775c4b8df;
			11'h3fe: dataout<=36'h7c9678aa8;
			11'h3ff: dataout<=36'h563368583;
			11'h400: dataout<=36'h48101a724;
			11'h401: dataout<=36'h771ccbb6c;
			11'h402: dataout<=36'h7cd1f8ea8;
			11'h403: dataout<=36'h5734a8937;
			11'h404: dataout<=36'h47c7da7e8;
			11'h405: dataout<=36'h76dc4bdf5;
			11'h406: dataout<=36'h7d0ab92a6;
			11'h407: dataout<=36'h5833a8cf6;
			11'h408: dataout<=36'h477f5a8ac;
			11'h409: dataout<=36'h769b0c07e;
			11'h40a: dataout<=36'h7d41f96a8;
			11'h40b: dataout<=36'h592fe90c0;
			11'h40c: dataout<=36'h4736da96f;
			11'h40d: dataout<=36'h76590c305;
			11'h40e: dataout<=36'h7d76f9aab;
			11'h40f: dataout<=36'h5a29a9494;
			11'h410: dataout<=36'h46eddaa31;
			11'h411: dataout<=36'h76158c58c;
			11'h412: dataout<=36'h7da979eb3;
			11'h413: dataout<=36'h5b20a9874;
			11'h414: dataout<=36'h46a51aaf3;
			11'h415: dataout<=36'h75d1cc811;
			11'h416: dataout<=36'h7ddaba2ba;
			11'h417: dataout<=36'h5c1529c5d;
			11'h418: dataout<=36'h465c1abb4;
			11'h419: dataout<=36'h758d4ca95;
			11'h41a: dataout<=36'h7e09ba6c3;
			11'h41b: dataout<=36'h5d06aa051;
			11'h41c: dataout<=36'h4612dac74;
			11'h41d: dataout<=36'h75474cd18;
			11'h41e: dataout<=36'h7e367aacf;
			11'h41f: dataout<=36'h5df5aa450;
			11'h420: dataout<=36'h45c99ad33;
			11'h421: dataout<=36'h7500ccf98;
			11'h422: dataout<=36'h7e60faeda;
			11'h423: dataout<=36'h5ee1ea858;
			11'h424: dataout<=36'h45805adf1;
			11'h425: dataout<=36'h74b98d216;
			11'h426: dataout<=36'h7e897b2e6;
			11'h427: dataout<=36'h5fcb6ac6b;
			11'h428: dataout<=36'h4536daeaf;
			11'h429: dataout<=36'h74718d494;
			11'h42a: dataout<=36'h7eb03b6f4;
			11'h42b: dataout<=36'h60b22b087;
			11'h42c: dataout<=36'h44ed1af6c;
			11'h42d: dataout<=36'h74284d710;
			11'h42e: dataout<=36'h7ed47bb05;
			11'h42f: dataout<=36'h6195eb4ad;
			11'h430: dataout<=36'h44a35b028;
			11'h431: dataout<=36'h73de8d98a;
			11'h432: dataout<=36'h7ef6fbf15;
			11'h433: dataout<=36'h6276eb8dd;
			11'h434: dataout<=36'h44595b0e3;
			11'h435: dataout<=36'h73938dc03;
			11'h436: dataout<=36'h7f16fc327;
			11'h437: dataout<=36'h63552bd17;
			11'h438: dataout<=36'h440f5b19d;
			11'h439: dataout<=36'h7347cde79;
			11'h43a: dataout<=36'h7f34bc739;
			11'h43b: dataout<=36'h64306c159;
			11'h43c: dataout<=36'h43c55b257;
			11'h43d: dataout<=36'h72fbce0ef;
			11'h43e: dataout<=36'h7f513cb4c;
			11'h43f: dataout<=36'h6508ac5a6;
			11'h440: dataout<=36'h437b1b310;
			11'h441: dataout<=36'h72ae8e363;
			11'h442: dataout<=36'h7f6b7cf61;
			11'h443: dataout<=36'h65ddec9fb;
			11'h444: dataout<=36'h43309b3c8;
			11'h445: dataout<=36'h72600e5d5;
			11'h446: dataout<=36'h7f82bd377;
			11'h447: dataout<=36'h66b06ce59;
			11'h448: dataout<=36'h42e61b47f;
			11'h449: dataout<=36'h72114e845;
			11'h44a: dataout<=36'h7f98bd78c;
			11'h44b: dataout<=36'h677fed2c1;
			11'h44c: dataout<=36'h429b5b536;
			11'h44d: dataout<=36'h71c14eab5;
			11'h44e: dataout<=36'h7fac7dba5;
			11'h44f: dataout<=36'h684c2d731;
			11'h450: dataout<=36'h42509b5eb;
			11'h451: dataout<=36'h71708ed21;
			11'h452: dataout<=36'h7fbd7dfbb;
			11'h453: dataout<=36'h69156dbaa;
			11'h454: dataout<=36'h4205db6a0;
			11'h455: dataout<=36'h711f4ef8c;
			11'h456: dataout<=36'h7fcd3e3d2;
			11'h457: dataout<=36'h69dbae02b;
			11'h458: dataout<=36'h41badb754;
			11'h459: dataout<=36'h70cd0f1f6;
			11'h45a: dataout<=36'h7fdabe7eb;
			11'h45b: dataout<=36'h6a9eee4b5;
			11'h45c: dataout<=36'h416f9b808;
			11'h45d: dataout<=36'h707a0f45f;
			11'h45e: dataout<=36'h7fe63ec05;
			11'h45f: dataout<=36'h6b5eee947;
			11'h460: dataout<=36'h41245b8ba;
			11'h461: dataout<=36'h7025cf6c4;
			11'h462: dataout<=36'h7feeff01d;
			11'h463: dataout<=36'h6c1beede1;
			11'h464: dataout<=36'h40d91b96c;
			11'h465: dataout<=36'h6fd18f929;
			11'h466: dataout<=36'h7ff6bf436;
			11'h467: dataout<=36'h6cd5af283;
			11'h468: dataout<=36'h408d9ba1d;
			11'h469: dataout<=36'h6f7bcfb8b;
			11'h46a: dataout<=36'h7ffb7f850;
			11'h46b: dataout<=36'h6d8c2f72d;
			11'h46c: dataout<=36'h40421bacd;
			11'h46d: dataout<=36'h6f25cfdec;
			11'h46e: dataout<=36'h7ffebfc69;
			11'h46f: dataout<=36'h6e3fafbde;
			11'h470: dataout<=36'h3ff65bb7c;
			11'h471: dataout<=36'h6ece5004a;
			11'h472: dataout<=36'h7fff00082;
			11'h473: dataout<=36'h6eefb0098;
			11'h474: dataout<=36'h3faa5bc2a;
			11'h475: dataout<=36'h6e76102a7;
			11'h476: dataout<=36'h7ffd4049d;
			11'h477: dataout<=36'h6f9cb0559;
			11'h478: dataout<=36'h3f5e9bcd8;
			11'h479: dataout<=36'h6e1d90502;
			11'h47a: dataout<=36'h7ffa408b6;
			11'h47b: dataout<=36'h704670a21;
			11'h47c: dataout<=36'h3f125bd85;
			11'h47d: dataout<=36'h6dc3d075c;
			11'h47e: dataout<=36'h7ff480cd1;
			11'h47f: dataout<=36'h70ecb0ef0;
			11'h480: dataout<=36'h3ec65be31;
			11'h481: dataout<=36'h6d69909b2;
			11'h482: dataout<=36'h7fed010e8;
			11'h483: dataout<=36'h718ff13c6;
			11'h484: dataout<=36'h3e79dbedc;
			11'h485: dataout<=36'h6d0e10c08;
			11'h486: dataout<=36'h7fe301503;
			11'h487: dataout<=36'h722fb18a3;
			11'h488: dataout<=36'h3e2d9bf87;
			11'h489: dataout<=36'h6cb290e5c;
			11'h48a: dataout<=36'h7fd80191b;
			11'h48b: dataout<=36'h72cc31d87;
			11'h48c: dataout<=36'h3de11c030;
			11'h48d: dataout<=36'h6c55910ac;
			11'h48e: dataout<=36'h7fc981d33;
			11'h48f: dataout<=36'h736532272;
			11'h490: dataout<=36'h3d945c0d9;
			11'h491: dataout<=36'h6bf7d12fc;
			11'h492: dataout<=36'h7fb98214c;
			11'h493: dataout<=36'h73faf2763;
			11'h494: dataout<=36'h3d479c181;
			11'h495: dataout<=36'h6b999154a;
			11'h496: dataout<=36'h7fa782563;
			11'h497: dataout<=36'h748d32c5a;
			11'h498: dataout<=36'h3cfadc228;
			11'h499: dataout<=36'h6b3a91794;
			11'h49a: dataout<=36'h7f9342978;
			11'h49b: dataout<=36'h751c33158;
			11'h49c: dataout<=36'h3caddc2ce;
			11'h49d: dataout<=36'h6ada919dd;
			11'h49e: dataout<=36'h7f7cc2d8e;
			11'h49f: dataout<=36'h75a7b365b;
			11'h4a0: dataout<=36'h3c60dc374;
			11'h4a1: dataout<=36'h6a7a11c25;
			11'h4a2: dataout<=36'h7f64c31a4;
			11'h4a3: dataout<=36'h762ff3b65;
			11'h4a4: dataout<=36'h3c139c418;
			11'h4a5: dataout<=36'h6a1851e69;
			11'h4a6: dataout<=36'h7f49c35b7;
			11'h4a7: dataout<=36'h76b474074;
			11'h4a8: dataout<=36'h3bc65c4bc;
			11'h4a9: dataout<=36'h69b6520ac;
			11'h4aa: dataout<=36'h7f2d839ca;
			11'h4ab: dataout<=36'h7735b4589;
			11'h4ac: dataout<=36'h3b78dc55f;
			11'h4ad: dataout<=36'h6953122ee;
			11'h4ae: dataout<=36'h7f0ec3dde;
			11'h4af: dataout<=36'h77b374aa3;
			11'h4b0: dataout<=36'h3b2b5c601;
			11'h4b1: dataout<=36'h68ef5252c;
			11'h4b2: dataout<=36'h7eee041ef;
			11'h4b3: dataout<=36'h782d74fc2;
			11'h4b4: dataout<=36'h3add9c6a3;
			11'h4b5: dataout<=36'h688a9276a;
			11'h4b6: dataout<=36'h7ecb04602;
			11'h4b7: dataout<=36'h78a4354e7;
			11'h4b8: dataout<=36'h3a901c743;
			11'h4b9: dataout<=36'h6825929a3;
			11'h4ba: dataout<=36'h7ea644a0e;
			11'h4bb: dataout<=36'h791775a11;
			11'h4bc: dataout<=36'h3a421c7e3;
			11'h4bd: dataout<=36'h67bf52bdd;
			11'h4be: dataout<=36'h7e7f44e1e;
			11'h4bf: dataout<=36'h7986f5f3f;
			11'h4c0: dataout<=36'h39f41c882;
			11'h4c1: dataout<=36'h675852e13;
			11'h4c2: dataout<=36'h7e564522c;
			11'h4c3: dataout<=36'h79f336472;
			11'h4c4: dataout<=36'h39a61c920;
			11'h4c5: dataout<=36'h66f0d3047;
			11'h4c6: dataout<=36'h7e2b05637;
			11'h4c7: dataout<=36'h7a5bb69aa;
			11'h4c8: dataout<=36'h39581c9bd;
			11'h4c9: dataout<=36'h6688d3278;
			11'h4ca: dataout<=36'h7dfe45a3f;
			11'h4cb: dataout<=36'h7ac0b6ee6;
			11'h4cc: dataout<=36'h3909dca59;
			11'h4cd: dataout<=36'h661f934a6;
			11'h4ce: dataout<=36'h7dce85e46;
			11'h4cf: dataout<=36'h7b21f7427;
			11'h4d0: dataout<=36'h38bb5caf5;
			11'h4d1: dataout<=36'h65b5936d5;
			11'h4d2: dataout<=36'h7d9d46250;
			11'h4d3: dataout<=36'h7b7fb796b;
			11'h4d4: dataout<=36'h386cdcb8f;
			11'h4d5: dataout<=36'h654ad38ff;
			11'h4d6: dataout<=36'h7d6986654;
			11'h4d7: dataout<=36'h7bd9f7eb3;
			11'h4d8: dataout<=36'h381e5cc29;
			11'h4d9: dataout<=36'h64df93b28;
			11'h4da: dataout<=36'h7d3406a58;
			11'h4db: dataout<=36'h7c3078400;
			11'h4dc: dataout<=36'h37cf9ccc2;
			11'h4dd: dataout<=36'h647353d4e;
			11'h4de: dataout<=36'h7cfc46e5a;
			11'h4df: dataout<=36'h7c837894f;
			11'h4e0: dataout<=36'h3780dcd5a;
			11'h4e1: dataout<=36'h640693f72;
			11'h4e2: dataout<=36'h7cc2c725a;
			11'h4e3: dataout<=36'h7cd2b8ea3;
			11'h4e4: dataout<=36'h37321cdf2;
			11'h4e5: dataout<=36'h639994195;
			11'h4e6: dataout<=36'h7c8807659;
			11'h4e7: dataout<=36'h7d1e793f9;
			11'h4e8: dataout<=36'h36e31ce88;
			11'h4e9: dataout<=36'h632b143b3;
			11'h4ea: dataout<=36'h7c49c7a54;
			11'h4eb: dataout<=36'h7d6679953;
			11'h4ec: dataout<=36'h3693dcf1e;
			11'h4ed: dataout<=36'h62bbd45d1;
			11'h4ee: dataout<=36'h7c09c7e50;
			11'h4ef: dataout<=36'h7daab9eaf;
			11'h4f0: dataout<=36'h3644dcfb3;
			11'h4f1: dataout<=36'h624c947ec;
			11'h4f2: dataout<=36'h7bc8c8248;
			11'h4f3: dataout<=36'h7deb7a40f;
			11'h4f4: dataout<=36'h35f59d046;
			11'h4f5: dataout<=36'h61dc14a02;
			11'h4f6: dataout<=36'h7b848863b;
			11'h4f7: dataout<=36'h7e287a971;
			11'h4f8: dataout<=36'h35a61d0da;
			11'h4f9: dataout<=36'h616ad4c1a;
			11'h4fa: dataout<=36'h7b3ec8a32;
			11'h4fb: dataout<=36'h7e61baed6;
			11'h4fc: dataout<=36'h35569d16c;
			11'h4fd: dataout<=36'h60f8d4e2d;
			11'h4fe: dataout<=36'h7af6c8e24;
			11'h4ff: dataout<=36'h7e977b43d;
			11'h500: dataout<=36'h35071d1fd;
			11'h501: dataout<=36'h60865503d;
			11'h502: dataout<=36'h7aacc9211;
			11'h503: dataout<=36'h7ec93b9a6;
			11'h504: dataout<=36'h34b75d28e;
			11'h505: dataout<=36'h60131524d;
			11'h506: dataout<=36'h7a6109600;
			11'h507: dataout<=36'h7ef77bf12;
			11'h508: dataout<=36'h34679d31d;
			11'h509: dataout<=36'h5f9f15458;
			11'h50a: dataout<=36'h7a13099e9;
			11'h50b: dataout<=36'h7f21fc47f;
			11'h50c: dataout<=36'h3417dd3ac;
			11'h50d: dataout<=36'h5f2a95661;
			11'h50e: dataout<=36'h79c349dd0;
			11'h50f: dataout<=36'h7f48bc9ee;
			11'h510: dataout<=36'h33c7dd43a;
			11'h511: dataout<=36'h5eb515868;
			11'h512: dataout<=36'h79714a1b6;
			11'h513: dataout<=36'h7f6bfcf5f;
			11'h514: dataout<=36'h3377dd4c7;
			11'h515: dataout<=36'h5e3f55a6d;
			11'h516: dataout<=36'h791d8a598;
			11'h517: dataout<=36'h7f8b3d4d1;
			11'h518: dataout<=36'h33279d554;
			11'h519: dataout<=36'h5dc855c70;
			11'h51a: dataout<=36'h78c78a97a;
			11'h51b: dataout<=36'h7fa6fda44;
			11'h51c: dataout<=36'h32d75d5df;
			11'h51d: dataout<=36'h5d50d5e6f;
			11'h51e: dataout<=36'h786f8ad57;
			11'h51f: dataout<=36'h7fbefdfb8;
			11'h520: dataout<=36'h32871d66a;
			11'h521: dataout<=36'h5cd91606d;
			11'h522: dataout<=36'h78164b132;
			11'h523: dataout<=36'h7fd2fe52d;
			11'h524: dataout<=36'h32369d6f3;
			11'h525: dataout<=36'h5c6016266;
			11'h526: dataout<=36'h77ba0b508;
			11'h527: dataout<=36'h7fe37eaa4;
			11'h528: dataout<=36'h31e61d77c;
			11'h529: dataout<=36'h5be69645e;
			11'h52a: dataout<=36'h775c0b8dd;
			11'h52b: dataout<=36'h7ff03f01a;
			11'h52c: dataout<=36'h31959d804;
			11'h52d: dataout<=36'h5b6c96653;
			11'h52e: dataout<=36'h76fc8bcae;
			11'h52f: dataout<=36'h7ff93f591;
			11'h530: dataout<=36'h3144dd88b;
			11'h531: dataout<=36'h5af1d6845;
			11'h532: dataout<=36'h769acc07b;
			11'h533: dataout<=36'h7ffe7fb09;
			11'h534: dataout<=36'h30f41d911;
			11'h535: dataout<=36'h5a7656a35;
			11'h536: dataout<=36'h76370c446;
			11'h537: dataout<=36'h7fffc0080;
			11'h538: dataout<=36'h30a35d997;
			11'h539: dataout<=36'h59fa96c23;
			11'h53a: dataout<=36'h75d20c80e;
			11'h53b: dataout<=36'h7ffdc05f7;
			11'h53c: dataout<=36'h30525da1b;
			11'h53d: dataout<=36'h597d96e0c;
			11'h53e: dataout<=36'h756a0cbd2;
			11'h53f: dataout<=36'h7ff7c0b6f;
			11'h540: dataout<=36'h30011da9f;
			11'h541: dataout<=36'h58ffd6ff6;
			11'h542: dataout<=36'h75008cf96;
			11'h543: dataout<=36'h7fee010e6;
			11'h544: dataout<=36'h2fb01db22;
			11'h545: dataout<=36'h5882171db;
			11'h546: dataout<=36'h74958d353;
			11'h547: dataout<=36'h7fe08165c;
			11'h548: dataout<=36'h2f5eddba4;
			11'h549: dataout<=36'h5803573be;
			11'h54a: dataout<=36'h74284d70e;
			11'h54b: dataout<=36'h7fcf81bd2;
			11'h54c: dataout<=36'h2f0d9dc25;
			11'h54d: dataout<=36'h57841759d;
			11'h54e: dataout<=36'h73b90dac4;
			11'h54f: dataout<=36'h7fba82147;
			11'h550: dataout<=36'h2ebc1dca5;
			11'h551: dataout<=36'h57041777a;
			11'h552: dataout<=36'h7347cde77;
			11'h553: dataout<=36'h7fa2026bc;
			11'h554: dataout<=36'h2e6a9dd24;
			11'h555: dataout<=36'h568357954;
			11'h556: dataout<=36'h72d48e226;
			11'h557: dataout<=36'h7f85c2c2f;
			11'h558: dataout<=36'h2e191dda3;
			11'h559: dataout<=36'h560257b2d;
			11'h55a: dataout<=36'h72604e5d3;
			11'h55b: dataout<=36'h7f65831a0;
			11'h55c: dataout<=36'h2dc75de20;
			11'h55d: dataout<=36'h558017d01;
			11'h55e: dataout<=36'h71e90e97b;
			11'h55f: dataout<=36'h7f41c3711;
			11'h560: dataout<=36'h2d75dde9d;
			11'h561: dataout<=36'h54fe17ed3;
			11'h562: dataout<=36'h71710ed1e;
			11'h563: dataout<=36'h7f1a43c7f;
			11'h564: dataout<=36'h2d23ddf19;
			11'h565: dataout<=36'h547a980a3;
			11'h566: dataout<=36'h70f64f0c0;
			11'h567: dataout<=36'h7eef041ec;
			11'h568: dataout<=36'h2cd21df94;
			11'h569: dataout<=36'h53f71826f;
			11'h56a: dataout<=36'h707a0f45c;
			11'h56b: dataout<=36'h7ec044757;
			11'h56c: dataout<=36'h2c801e00e;
			11'h56d: dataout<=36'h5372d8438;
			11'h56e: dataout<=36'h6ffc0f7f3;
			11'h56f: dataout<=36'h7e8d84cc0;
			11'h570: dataout<=36'h2c2e1e087;
			11'h571: dataout<=36'h52edd85ff;
			11'h572: dataout<=36'h6f7c0fb87;
			11'h573: dataout<=36'h7e5745227;
			11'h574: dataout<=36'h2bdbde100;
			11'h575: dataout<=36'h5268187c4;
			11'h576: dataout<=36'h6efa0ff1a;
			11'h577: dataout<=36'h7e1d4578b;
			11'h578: dataout<=36'h2b899e177;
			11'h579: dataout<=36'h51e1d8984;
			11'h57a: dataout<=36'h6e76102a4;
			11'h57b: dataout<=36'h7ddfc5ced;
			11'h57c: dataout<=36'h2b375e1ee;
			11'h57d: dataout<=36'h515b58b43;
			11'h57e: dataout<=36'h6df11062d;
			11'h57f: dataout<=36'h7d9e4624c;
			11'h580: dataout<=36'h2ae4de263;
			11'h581: dataout<=36'h50d398cfe;
			11'h582: dataout<=36'h6d69509b0;
			11'h583: dataout<=36'h7d59467a8;
			11'h584: dataout<=36'h2a925e2d8;
			11'h585: dataout<=36'h504b98eb7;
			11'h586: dataout<=36'h6ce010d30;
			11'h587: dataout<=36'h7d1086d01;
			11'h588: dataout<=36'h2a3fde34c;
			11'h589: dataout<=36'h4fc31906c;
			11'h58a: dataout<=36'h6c55510aa;
			11'h58b: dataout<=36'h7cc447257;
			11'h58c: dataout<=36'h29ed5e3bf;
			11'h58d: dataout<=36'h4f3a1921e;
			11'h58e: dataout<=36'h6bc8d141f;
			11'h58f: dataout<=36'h7c74477aa;
			11'h590: dataout<=36'h299a9e431;
			11'h591: dataout<=36'h4eb0593ce;
			11'h592: dataout<=36'h6b3a51791;
			11'h593: dataout<=36'h7c20c7cf9;
			11'h594: dataout<=36'h2947de4a3;
			11'h595: dataout<=36'h4e265957c;
			11'h596: dataout<=36'h6aaa91b00;
			11'h597: dataout<=36'h7bc988244;
			11'h598: dataout<=36'h28f51e513;
			11'h599: dataout<=36'h4d9b99725;
			11'h59a: dataout<=36'h6a1891e67;
			11'h59b: dataout<=36'h7b6ec878c;
			11'h59c: dataout<=36'h28a21e583;
			11'h59d: dataout<=36'h4d10198cd;
			11'h59e: dataout<=36'h6985121cc;
			11'h59f: dataout<=36'h7b1048cd0;
			11'h5a0: dataout<=36'h284f1e5f1;
			11'h5a1: dataout<=36'h4c83d9a6f;
			11'h5a2: dataout<=36'h68ef12529;
			11'h5a3: dataout<=36'h7aae4920f;
			11'h5a4: dataout<=36'h27fc1e65f;
			11'h5a5: dataout<=36'h4bf799c11;
			11'h5a6: dataout<=36'h685852884;
			11'h5a7: dataout<=36'h7a488974b;
			11'h5a8: dataout<=36'h27a8de6cc;
			11'h5a9: dataout<=36'h4b6a59daf;
			11'h5aa: dataout<=36'h67bf52bda;
			11'h5ab: dataout<=36'h79df89c81;
			11'h5ac: dataout<=36'h27559e738;
			11'h5ad: dataout<=36'h4adc99f4a;
			11'h5ae: dataout<=36'h6724d2f2b;
			11'h5af: dataout<=36'h7972ca1b4;
			11'h5b0: dataout<=36'h27025e7a3;
			11'h5b1: dataout<=36'h4a4e5a0e1;
			11'h5b2: dataout<=36'h668853276;
			11'h5b3: dataout<=36'h79028a6e1;
			11'h5b4: dataout<=36'h26af1e80d;
			11'h5b5: dataout<=36'h49bfda276;
			11'h5b6: dataout<=36'h65ead35bc;
			11'h5b7: dataout<=36'h788e8ac0a;
			11'h5b8: dataout<=36'h265b9e876;
			11'h5b9: dataout<=36'h49305a407;
			11'h5ba: dataout<=36'h654ad38fd;
			11'h5bb: dataout<=36'h78174b12e;
			11'h5bc: dataout<=36'h26081e8df;
			11'h5bd: dataout<=36'h48a09a597;
			11'h5be: dataout<=36'h64a9d3c3b;
			11'h5bf: dataout<=36'h779c8b64c;
			11'h5c0: dataout<=36'h25b49e946;
			11'h5c1: dataout<=36'h48105a721;
			11'h5c2: dataout<=36'h6406d3f6f;
			11'h5c3: dataout<=36'h771e0bb66;
			11'h5c4: dataout<=36'h2560de9ad;
			11'h5c5: dataout<=36'h477f5a8aa;
			11'h5c6: dataout<=36'h6362142a2;
			11'h5c7: dataout<=36'h769c4c079;
			11'h5c8: dataout<=36'h250d5ea13;
			11'h5c9: dataout<=36'h46ee5aa30;
			11'h5ca: dataout<=36'h62bc545cf;
			11'h5cb: dataout<=36'h76170c588;
			11'h5cc: dataout<=36'h24b99ea78;
			11'h5cd: dataout<=36'h465c9abb2;
			11'h5ce: dataout<=36'h6214d48f5;
			11'h5cf: dataout<=36'h758e4ca90;
			11'h5d0: dataout<=36'h24659eadb;
			11'h5d1: dataout<=36'h45c99ad30;
			11'h5d2: dataout<=36'h616a54c16;
			11'h5d3: dataout<=36'h75024cf92;
			11'h5d4: dataout<=36'h2411deb3f;
			11'h5d5: dataout<=36'h45371aeae;
			11'h5d6: dataout<=36'h60c054f34;
			11'h5d7: dataout<=36'h74728d48f;
			11'h5d8: dataout<=36'h23bddeba1;
			11'h5d9: dataout<=36'h44a39b026;
			11'h5da: dataout<=36'h60135524a;
			11'h5db: dataout<=36'h73df8d985;
			11'h5dc: dataout<=36'h2369dec02;
			11'h5dd: dataout<=36'h440fdb19b;
			11'h5de: dataout<=36'h5f655555a;
			11'h5df: dataout<=36'h73494de75;
			11'h5e0: dataout<=36'h23159ec62;
			11'h5e1: dataout<=36'h437b1b30e;
			11'h5e2: dataout<=36'h5eb515867;
			11'h5e3: dataout<=36'h72af8e35e;
			11'h5e4: dataout<=36'h22c19ecc2;
			11'h5e5: dataout<=36'h42e69b47e;
			11'h5e6: dataout<=36'h5e0495b6d;
			11'h5e7: dataout<=36'h72128e841;
			11'h5e8: dataout<=36'h226d5ed20;
			11'h5e9: dataout<=36'h42511b5e9;
			11'h5ea: dataout<=36'h5d5155e6c;
			11'h5eb: dataout<=36'h71720ed1d;
			11'h5ec: dataout<=36'h22191ed7e;
			11'h5ed: dataout<=36'h41bb1b752;
			11'h5ee: dataout<=36'h5c9cd6166;
			11'h5ef: dataout<=36'h70ce8f1f2;
			11'h5f0: dataout<=36'h21c49eddb;
			11'h5f1: dataout<=36'h41249b8b9;
			11'h5f2: dataout<=36'h5be6d645d;
			11'h5f3: dataout<=36'h70278f6c0;
			11'h5f4: dataout<=36'h21705ee37;
			11'h5f5: dataout<=36'h408e1ba1b;
			11'h5f6: dataout<=36'h5b2fd674b;
			11'h5f7: dataout<=36'h6f7d4fb87;
			11'h5f8: dataout<=36'h211bdee92;
			11'h5f9: dataout<=36'h3ff69bb7b;
			11'h5fa: dataout<=36'h5a76d6a34;
			11'h5fb: dataout<=36'h6ecf90046;
			11'h5fc: dataout<=36'h20c75eeec;
			11'h5fd: dataout<=36'h3f5f1bcd7;
			11'h5fe: dataout<=36'h59bcd6d17;
			11'h5ff: dataout<=36'h6e1ed04fe;
			11'h600: dataout<=36'h20729ef45;
			11'h601: dataout<=36'h3ec65be30;
			11'h602: dataout<=36'h590016ff5;
			11'h603: dataout<=36'h6d6b109ae;
			11'h604: dataout<=36'h201e1ef9d;
			11'h605: dataout<=36'h3e2e1bf84;
			11'h606: dataout<=36'h5843572c9;
			11'h607: dataout<=36'h6cb3d0e57;
			11'h608: dataout<=36'h1fc95eff4;
			11'h609: dataout<=36'h3d949c0d6;
			11'h60a: dataout<=36'h57841759a;
			11'h60b: dataout<=36'h6bf9912f7;
			11'h60c: dataout<=36'h1f749f04b;
			11'h60d: dataout<=36'h3cfb1c226;
			11'h60e: dataout<=36'h56c417865;
			11'h60f: dataout<=36'h6b3c11790;
			11'h610: dataout<=36'h1f1f9f0a0;
			11'h611: dataout<=36'h3c60dc371;
			11'h612: dataout<=36'h560217b29;
			11'h613: dataout<=36'h6a7b51c21;
			11'h614: dataout<=36'h1ecadf0f5;
			11'h615: dataout<=36'h3bc69c4ba;
			11'h616: dataout<=36'h553f57de8;
			11'h617: dataout<=36'h69b7920a9;
			11'h618: dataout<=36'h1e75df149;
			11'h619: dataout<=36'h3b2b9c600;
			11'h61a: dataout<=36'h547ad80a1;
			11'h61b: dataout<=36'h68f0d2528;
			11'h61c: dataout<=36'h1e20df19c;
			11'h61d: dataout<=36'h3a901c742;
			11'h61e: dataout<=36'h53b4d8353;
			11'h61f: dataout<=36'h6826d29a0;
			11'h620: dataout<=36'h1dcbdf1ed;
			11'h621: dataout<=36'h39f45c87f;
			11'h622: dataout<=36'h52ed985fc;
			11'h623: dataout<=36'h675a12e0e;
			11'h624: dataout<=36'h1d76df23e;
			11'h625: dataout<=36'h39585c9ba;
			11'h626: dataout<=36'h5225588a1;
			11'h627: dataout<=36'h668a13274;
			11'h628: dataout<=36'h1d219f28f;
			11'h629: dataout<=36'h38bb9caf4;
			11'h62a: dataout<=36'h515b58b42;
			11'h62b: dataout<=36'h65b7136d1;
			11'h62c: dataout<=36'h1ccc5f2de;
			11'h62d: dataout<=36'h381e9cc28;
			11'h62e: dataout<=36'h509018dda;
			11'h62f: dataout<=36'h64e153b24;
			11'h630: dataout<=36'h1c771f32c;
			11'h631: dataout<=36'h37811cd59;
			11'h632: dataout<=36'h4fc35906b;
			11'h633: dataout<=36'h640853f6f;
			11'h634: dataout<=36'h1c21df379;
			11'h635: dataout<=36'h36e35ce86;
			11'h636: dataout<=36'h4ef5992f4;
			11'h637: dataout<=36'h632c943b0;
			11'h638: dataout<=36'h1bcc5f3c6;
			11'h639: dataout<=36'h3644dcfb1;
			11'h63a: dataout<=36'h4e261957a;
			11'h63b: dataout<=36'h624e147e8;
			11'h63c: dataout<=36'h1b771f411;
			11'h63d: dataout<=36'h35a69d0d7;
			11'h63e: dataout<=36'h4d56197f5;
			11'h63f: dataout<=36'h616c54c16;
			11'h640: dataout<=36'h1b219f45c;
			11'h641: dataout<=36'h35075d1fb;
			11'h642: dataout<=36'h4c8419a6d;
			11'h643: dataout<=36'h60881503a;
			11'h644: dataout<=36'h1acc1f4a6;
			11'h645: dataout<=36'h34681d31c;
			11'h646: dataout<=36'h4bb159cde;
			11'h647: dataout<=36'h5fa0d5455;
			11'h648: dataout<=36'h1a769f4ef;
			11'h649: dataout<=36'h33c85d439;
			11'h64a: dataout<=36'h4add59f48;
			11'h64b: dataout<=36'h5eb6d5866;
			11'h64c: dataout<=36'h1a20df536;
			11'h64d: dataout<=36'h3327dd551;
			11'h64e: dataout<=36'h4a075a1a9;
			11'h64f: dataout<=36'h5dca15c6c;
			11'h650: dataout<=36'h19cb5f57d;
			11'h651: dataout<=36'h32879d667;
			11'h652: dataout<=36'h49311a404;
			11'h653: dataout<=36'h5cda96069;
			11'h654: dataout<=36'h19759f5c3;
			11'h655: dataout<=36'h31e69d779;
			11'h656: dataout<=36'h4858da658;
			11'h657: dataout<=36'h5be89645b;
			11'h658: dataout<=36'h191fdf609;
			11'h659: dataout<=36'h31455d88a;
			11'h65a: dataout<=36'h47801a8a9;
			11'h65b: dataout<=36'h5af396843;
			11'h65c: dataout<=36'h18ca1f64d;
			11'h65d: dataout<=36'h30a3dd995;
			11'h65e: dataout<=36'h46a61aaef;
			11'h65f: dataout<=36'h59fc16c20;
			11'h660: dataout<=36'h18741f690;
			11'h661: dataout<=36'h30019da9d;
			11'h662: dataout<=36'h45ca1ad2e;
			11'h663: dataout<=36'h5901d6ff2;
			11'h664: dataout<=36'h181e5f6d3;
			11'h665: dataout<=36'h2f5f5dba3;
			11'h666: dataout<=36'h44eddaf69;
			11'h667: dataout<=36'h5805173ba;
			11'h668: dataout<=36'h17c85f714;
			11'h669: dataout<=36'h2ebc9dca3;
			11'h66a: dataout<=36'h44101b199;
			11'h66b: dataout<=36'h5705d7777;
			11'h66c: dataout<=36'h17725f755;
			11'h66d: dataout<=36'h2e199dda2;
			11'h66e: dataout<=36'h43315b3c5;
			11'h66f: dataout<=36'h5603d7b29;
			11'h670: dataout<=36'h171c5f794;
			11'h671: dataout<=36'h2d761de9b;
			11'h672: dataout<=36'h42515b5e7;
			11'h673: dataout<=36'h54ff97ed0;
			11'h674: dataout<=36'h16c65f7d3;
			11'h675: dataout<=36'h2cd29df92;
			11'h676: dataout<=36'h41709b803;
			11'h677: dataout<=36'h53f8d826c;
			11'h678: dataout<=36'h16701f811;
			11'h679: dataout<=36'h2c2e5e086;
			11'h67a: dataout<=36'h408e1ba1a;
			11'h67b: dataout<=36'h52ef585fd;
			11'h67c: dataout<=36'h161a1f84e;
			11'h67d: dataout<=36'h2b8a1e176;
			11'h67e: dataout<=36'h3fab5bc27;
			11'h67f: dataout<=36'h51e398982;
			11'h680: dataout<=36'h15c3df88a;
			11'h681: dataout<=36'h2ae55e263;
			11'h682: dataout<=36'h3ec71be2f;
			11'h683: dataout<=36'h50d598cfc;
			11'h684: dataout<=36'h156d9f8c5;
			11'h685: dataout<=36'h2a405e34b;
			11'h686: dataout<=36'h3de1dc02d;
			11'h687: dataout<=36'h4fc51906a;
			11'h688: dataout<=36'h15175f8ff;
			11'h689: dataout<=36'h299b1e430;
			11'h68a: dataout<=36'h3cfb9c225;
			11'h68b: dataout<=36'h4eb2593cc;
			11'h68c: dataout<=36'h14c11f938;
			11'h68d: dataout<=36'h28f59e512;
			11'h68e: dataout<=36'h3c145c415;
			11'h68f: dataout<=36'h4d9d19723;
			11'h690: dataout<=36'h146a9f970;
			11'h691: dataout<=36'h284f5e5ef;
			11'h692: dataout<=36'h3b2b9c5fd;
			11'h693: dataout<=36'h4c85d9a6d;
			11'h694: dataout<=36'h14145f9a8;
			11'h695: dataout<=36'h27a95e6cb;
			11'h696: dataout<=36'h3a42dc7e0;
			11'h697: dataout<=36'h4b6c19dac;
			11'h698: dataout<=36'h13bddf9de;
			11'h699: dataout<=36'h27029e7a1;
			11'h69a: dataout<=36'h39585c9b9;
			11'h69b: dataout<=36'h4a505a0df;
			11'h69c: dataout<=36'h13675fa13;
			11'h69d: dataout<=36'h265bde874;
			11'h69e: dataout<=36'h386d1cb8b;
			11'h69f: dataout<=36'h49325a405;
			11'h6a0: dataout<=36'h13111fa48;
			11'h6a1: dataout<=36'h25b51e944;
			11'h6a2: dataout<=36'h3781dcd56;
			11'h6a3: dataout<=36'h48125a720;
			11'h6a4: dataout<=36'h12ba5fa7c;
			11'h6a5: dataout<=36'h250d5ea12;
			11'h6a6: dataout<=36'h36945cf1c;
			11'h6a7: dataout<=36'h46f01aa2e;
			11'h6a8: dataout<=36'h1263dfaae;
			11'h6a9: dataout<=36'h2465dead9;
			11'h6aa: dataout<=36'h35a65d0d5;
			11'h6ab: dataout<=36'h45cbdad2f;
			11'h6ac: dataout<=36'h120d5fae0;
			11'h6ad: dataout<=36'h23be5eb9f;
			11'h6ae: dataout<=36'h34b85d28a;
			11'h6af: dataout<=36'h44a55b024;
			11'h6b0: dataout<=36'h11b69fb11;
			11'h6b1: dataout<=36'h2315dec61;
			11'h6b2: dataout<=36'h33c81d437;
			11'h6b3: dataout<=36'h437d1b30c;
			11'h6b4: dataout<=36'h11601fb41;
			11'h6b5: dataout<=36'h226dded1e;
			11'h6b6: dataout<=36'h32d85d5da;
			11'h6b7: dataout<=36'h4252db5e8;
			11'h6b8: dataout<=36'h11095fb70;
			11'h6b9: dataout<=36'h21c51edd9;
			11'h6ba: dataout<=36'h31e6dd778;
			11'h6bb: dataout<=36'h41269b8b7;
			11'h6bc: dataout<=36'h10b29fb9e;
			11'h6bd: dataout<=36'h211c1ee90;
			11'h6be: dataout<=36'h30f49d90e;
			11'h6bf: dataout<=36'h3ff85bb79;
			11'h6c0: dataout<=36'h105bdfbcb;
			11'h6c1: dataout<=36'h2072def42;
			11'h6c2: dataout<=36'h30019da9a;
			11'h6c3: dataout<=36'h3ec85be2e;
			11'h6c4: dataout<=36'h10051fbf8;
			11'h6c5: dataout<=36'h1fc99eff3;
			11'h6c6: dataout<=36'h2f0e1dc22;
			11'h6c7: dataout<=36'h3d969c0d6;
			11'h6c8: dataout<=36'h0fae5fc23;
			11'h6c9: dataout<=36'h1f201f09f;
			11'h6ca: dataout<=36'h2e19ddd9f;
			11'h6cb: dataout<=36'h3c62dc370;
			11'h6cc: dataout<=36'h0f579fc4d;
			11'h6cd: dataout<=36'h1e769f146;
			11'h6ce: dataout<=36'h2d24ddf14;
			11'h6cf: dataout<=36'h3b2d9c5fe;
			11'h6d0: dataout<=36'h0f009fc77;
			11'h6d1: dataout<=36'h1dcc1f1ec;
			11'h6d2: dataout<=36'h2c2e9e084;
			11'h6d3: dataout<=36'h39f65c87f;
			11'h6d4: dataout<=36'h0ea9dfca0;
			11'h6d5: dataout<=36'h1d225f28e;
			11'h6d6: dataout<=36'h2b389e1eb;
			11'h6d7: dataout<=36'h38bd9caf2;
			11'h6d8: dataout<=36'h0e52dfcc7;
			11'h6d9: dataout<=36'h1c779f32a;
			11'h6da: dataout<=36'h2a40de348;
			11'h6db: dataout<=36'h37831cd58;
			11'h6dc: dataout<=36'h0dfbdfcee;
			11'h6dd: dataout<=36'h1bccdf3c5;
			11'h6de: dataout<=36'h29489e4a0;
			11'h6df: dataout<=36'h36471cfb0;
			11'h6e0: dataout<=36'h0da4dfd14;
			11'h6e1: dataout<=36'h1b21df45b;
			11'h6e2: dataout<=36'h284f9e5ef;
			11'h6e3: dataout<=36'h35095d1fb;
			11'h6e4: dataout<=36'h0d4ddfd38;
			11'h6e5: dataout<=36'h1a76df4ec;
			11'h6e6: dataout<=36'h27565e733;
			11'h6e7: dataout<=36'h33ca1d438;
			11'h6e8: dataout<=36'h0cf6dfd5c;
			11'h6e9: dataout<=36'h19cb9f57b;
			11'h6ea: dataout<=36'h265c5e872;
			11'h6eb: dataout<=36'h32895d667;
			11'h6ec: dataout<=36'h0c9fdfd7f;
			11'h6ed: dataout<=36'h19201f607;
			11'h6ee: dataout<=36'h25619e9a9;
			11'h6ef: dataout<=36'h31471d889;
			11'h6f0: dataout<=36'h0c48dfda1;
			11'h6f1: dataout<=36'h18749f68e;
			11'h6f2: dataout<=36'h24669ead7;
			11'h6f3: dataout<=36'h30039da9d;
			11'h6f4: dataout<=36'h0bf19fdc2;
			11'h6f5: dataout<=36'h17c85f712;
			11'h6f6: dataout<=36'h236a1ebfe;
			11'h6f7: dataout<=36'h2ebe5dca3;
			11'h6f8: dataout<=36'h0b9a9fde3;
			11'h6f9: dataout<=36'h171cdf794;
			11'h6fa: dataout<=36'h226e5ed1f;
			11'h6fb: dataout<=36'h2d781de9b;
			11'h6fc: dataout<=36'h0b439fe02;
			11'h6fd: dataout<=36'h1670df80f;
			11'h6fe: dataout<=36'h21715ee33;
			11'h6ff: dataout<=36'h2c305e085;
			11'h700: dataout<=36'h0aec5fe20;
			11'h701: dataout<=36'h15c45f888;
			11'h702: dataout<=36'h20739ef41;
			11'h703: dataout<=36'h2ae75e261;
			11'h704: dataout<=36'h0a951fe3e;
			11'h705: dataout<=36'h15179f8fe;
			11'h706: dataout<=36'h1f751f049;
			11'h707: dataout<=36'h299cde42f;
			11'h708: dataout<=36'h0a3e1fe5a;
			11'h709: dataout<=36'h146b5f96f;
			11'h70a: dataout<=36'h1e771f146;
			11'h70b: dataout<=36'h28515e5ef;
			11'h70c: dataout<=36'h09e6dfe76;
			11'h70d: dataout<=36'h13be9f9dd;
			11'h70e: dataout<=36'h1d77df23c;
			11'h70f: dataout<=36'h2704de7a1;
			11'h710: dataout<=36'h098f9fe90;
			11'h711: dataout<=36'h13119fa46;
			11'h712: dataout<=36'h1c781f328;
			11'h713: dataout<=36'h25b6de945;
			11'h714: dataout<=36'h09385feaa;
			11'h715: dataout<=36'h12645faad;
			11'h716: dataout<=36'h1b77df40e;
			11'h717: dataout<=36'h24681eada;
			11'h718: dataout<=36'h08e11fec3;
			11'h719: dataout<=36'h11b75fb11;
			11'h71a: dataout<=36'h1a779f4ed;
			11'h71b: dataout<=36'h23181ec61;
			11'h71c: dataout<=36'h0889dfeda;
			11'h71d: dataout<=36'h1109dfb6e;
			11'h71e: dataout<=36'h19765f5bf;
			11'h71f: dataout<=36'h21c71edd9;
			11'h720: dataout<=36'h08329fef1;
			11'h721: dataout<=36'h105c9fbc9;
			11'h722: dataout<=36'h18755f68c;
			11'h723: dataout<=36'h20751ef44;
			11'h724: dataout<=36'h07db1ff07;
			11'h725: dataout<=36'h0fae9fc21;
			11'h726: dataout<=36'h1772df751;
			11'h727: dataout<=36'h1f221f09f;
			11'h728: dataout<=36'h0783dff1c;
			11'h729: dataout<=36'h0f011fc75;
			11'h72a: dataout<=36'h16711f80d;
			11'h72b: dataout<=36'h1dce5f1ec;
			11'h72c: dataout<=36'h072c9ff30;
			11'h72d: dataout<=36'h0e535fcc5;
			11'h72e: dataout<=36'h156e9f8c1;
			11'h72f: dataout<=36'h1c799f32b;
			11'h730: dataout<=36'h06d51ff44;
			11'h731: dataout<=36'h0da51fd13;
			11'h732: dataout<=36'h146b5f96f;
			11'h733: dataout<=36'h1b241f45b;
			11'h734: dataout<=36'h067ddff56;
			11'h735: dataout<=36'h0cf75fd5c;
			11'h736: dataout<=36'h13685fa12;
			11'h737: dataout<=36'h19cd9f57d;
			11'h738: dataout<=36'h06265ff67;
			11'h739: dataout<=36'h0c491fda0;
			11'h73a: dataout<=36'h12649faac;
			11'h73b: dataout<=36'h18769f68f;
			11'h73c: dataout<=36'h05cf1ff77;
			11'h73d: dataout<=36'h0b9b1fde1;
			11'h73e: dataout<=36'h11611fb3e;
			11'h73f: dataout<=36'h171edf794;
			11'h740: dataout<=36'h05779ff87;
			11'h741: dataout<=36'h0aec9fe1f;
			11'h742: dataout<=36'h105c9fbc9;
			11'h743: dataout<=36'h15c65f889;
			11'h744: dataout<=36'h05205ff95;
			11'h745: dataout<=36'h0a3e9fe58;
			11'h746: dataout<=36'h0f589fc4a;
			11'h747: dataout<=36'h146d1f970;
			11'h748: dataout<=36'h04c8dffa3;
			11'h749: dataout<=36'h09901fe8f;
			11'h74a: dataout<=36'h0e53dfcc5;
			11'h74b: dataout<=36'h13135fa48;
			11'h74c: dataout<=36'h04715ffaf;
			11'h74d: dataout<=36'h08e15fec1;
			11'h74e: dataout<=36'h0d4e9fd35;
			11'h74f: dataout<=36'h11b91fb11;
			11'h750: dataout<=36'h041a1ffbb;
			11'h751: dataout<=36'h08331fef0;
			11'h752: dataout<=36'h0c49dfd9f;
			11'h753: dataout<=36'h105e5fbcb;
			11'h754: dataout<=36'h03c29ffc6;
			11'h755: dataout<=36'h07845ff1b;
			11'h756: dataout<=36'h0b445fdff;
			11'h757: dataout<=36'h0f031fc77;
			11'h758: dataout<=36'h036b1ffd0;
			11'h759: dataout<=36'h06d59ff43;
			11'h75a: dataout<=36'h0a3edfe59;
			11'h75b: dataout<=36'h0da75fd14;
			11'h75c: dataout<=36'h03139ffd9;
			11'h75d: dataout<=36'h0626dff67;
			11'h75e: dataout<=36'h09391fea9;
			11'h75f: dataout<=36'h0c4b5fda2;
			11'h760: dataout<=36'h02bc5ffe1;
			11'h761: dataout<=36'h05785ff87;
			11'h762: dataout<=36'h0833dfef1;
			11'h763: dataout<=36'h0aeedfe21;
			11'h764: dataout<=36'h0264dffe8;
			11'h765: dataout<=36'h04c99ffa3;
			11'h766: dataout<=36'h072ddff30;
			11'h767: dataout<=36'h09921fe91;
			11'h768: dataout<=36'h020d5ffee;
			11'h769: dataout<=36'h041a9ffbb;
			11'h76a: dataout<=36'h06279ff66;
			11'h76b: dataout<=36'h0834dfef2;
			11'h76c: dataout<=36'h01b5dfff3;
			11'h76d: dataout<=36'h036b9ffcf;
			11'h76e: dataout<=36'h05215ff94;
			11'h76f: dataout<=36'h06d79ff44;
			11'h770: dataout<=36'h015e5fff7;
			11'h771: dataout<=36'h02bc9ffe0;
			11'h772: dataout<=36'h041adffba;
			11'h773: dataout<=36'h057a1ff87;
			11'h774: dataout<=36'h0106dfffa;
			11'h775: dataout<=36'h020d9ffec;
			11'h776: dataout<=36'h03145ffd6;
			11'h777: dataout<=36'h041c5ffbc;
			11'h778: dataout<=36'h00af5fffd;
			11'h779: dataout<=36'h015e9fff7;
			11'h77a: dataout<=36'h020ddffed;
			11'h77b: dataout<=36'h02be9ffe1;
			11'h77c: dataout<=36'h00af5fffd;
			11'h77d: dataout<=36'h015e9fff7;
			11'h77e: dataout<=36'h020ddffed;
			11'h77f: dataout<=36'h02be9ffe1;
			11'h780: dataout<=36'h000000000;
			11'h781: dataout<=36'h000000000;
			11'h782: dataout<=36'h000000000;
			11'h783: dataout<=36'h000000000;
			11'h784: dataout<=36'h000000000;
			11'h785: dataout<=36'h000000000;
			11'h786: dataout<=36'h000000000;
			11'h787: dataout<=36'h000000000;
			11'h788: dataout<=36'h000000000;
			11'h789: dataout<=36'h000000000;
			11'h78a: dataout<=36'h000000000;
			11'h78b: dataout<=36'h000000000;
			11'h78c: dataout<=36'h000000000;
			11'h78d: dataout<=36'h000000000;
			11'h78e: dataout<=36'h000000000;
			11'h78f: dataout<=36'h000000000;
			11'h790: dataout<=36'h000000000;
			11'h791: dataout<=36'h000000000;
			11'h792: dataout<=36'h000000000;
			11'h793: dataout<=36'h000000000;
			11'h794: dataout<=36'h000000000;
			11'h795: dataout<=36'h000000000;
			11'h796: dataout<=36'h000000000;
			11'h797: dataout<=36'h000000000;
			11'h798: dataout<=36'h000000000;
			11'h799: dataout<=36'h000000000;
			11'h79a: dataout<=36'h000000000;
			11'h79b: dataout<=36'h000000000;
			11'h79c: dataout<=36'h000000000;
			11'h79d: dataout<=36'h000000000;
			11'h79e: dataout<=36'h000000000;
			11'h79f: dataout<=36'h000000000;
			11'h7a0: dataout<=36'h000000000;
			11'h7a1: dataout<=36'h000000000;
			11'h7a2: dataout<=36'h000000000;
			11'h7a3: dataout<=36'h000000000;
			11'h7a4: dataout<=36'h000000000;
			11'h7a5: dataout<=36'h000000000;
			11'h7a6: dataout<=36'h000000000;
			11'h7a7: dataout<=36'h000000000;
			11'h7a8: dataout<=36'h000000000;
			11'h7a9: dataout<=36'h000000000;
			11'h7aa: dataout<=36'h000000000;
			11'h7ab: dataout<=36'h000000000;
			11'h7ac: dataout<=36'h000000000;
			11'h7ad: dataout<=36'h000000000;
			11'h7ae: dataout<=36'h000000000;
			11'h7af: dataout<=36'h000000000;
			11'h7b0: dataout<=36'h000000000;
			11'h7b1: dataout<=36'h000000000;
			11'h7b2: dataout<=36'h000000000;
			11'h7b3: dataout<=36'h000000000;
			11'h7b4: dataout<=36'h000000000;
			11'h7b5: dataout<=36'h000000000;
			11'h7b6: dataout<=36'h000000000;
			11'h7b7: dataout<=36'h000000000;
			11'h7b8: dataout<=36'h000000000;
			11'h7b9: dataout<=36'h000000000;
			11'h7ba: dataout<=36'h000000000;
			11'h7bb: dataout<=36'h000000000;
			11'h7bc: dataout<=36'h000000000;
			11'h7bd: dataout<=36'h000000000;
			11'h7be: dataout<=36'h000000000;
			11'h7bf: dataout<=36'h000000000;
			11'h7c0: dataout<=36'h000000000;
			11'h7c1: dataout<=36'h000000000;
			11'h7c2: dataout<=36'h000000000;
			11'h7c3: dataout<=36'h000000000;
			11'h7c4: dataout<=36'h000000000;
			11'h7c5: dataout<=36'h000000000;
			11'h7c6: dataout<=36'h000000000;
			11'h7c7: dataout<=36'h000000000;
			11'h7c8: dataout<=36'h000000000;
			11'h7c9: dataout<=36'h000000000;
			11'h7ca: dataout<=36'h000000000;
			11'h7cb: dataout<=36'h000000000;
			11'h7cc: dataout<=36'h000000000;
			11'h7cd: dataout<=36'h000000000;
			11'h7ce: dataout<=36'h000000000;
			11'h7cf: dataout<=36'h000000000;
			11'h7d0: dataout<=36'h000000000;
			11'h7d1: dataout<=36'h000000000;
			11'h7d2: dataout<=36'h000000000;
			11'h7d3: dataout<=36'h000000000;
			11'h7d4: dataout<=36'h000000000;
			11'h7d5: dataout<=36'h000000000;
			11'h7d6: dataout<=36'h000000000;
			11'h7d7: dataout<=36'h000000000;
			11'h7d8: dataout<=36'h000000000;
			11'h7d9: dataout<=36'h000000000;
			11'h7da: dataout<=36'h000000000;
			11'h7db: dataout<=36'h000000000;
			11'h7dc: dataout<=36'h000000000;
			11'h7dd: dataout<=36'h000000000;
			11'h7de: dataout<=36'h000000000;
			11'h7df: dataout<=36'h000000000;
			11'h7e0: dataout<=36'h000000000;
			11'h7e1: dataout<=36'h000000000;
			11'h7e2: dataout<=36'h000000000;
			11'h7e3: dataout<=36'h000000000;
			11'h7e4: dataout<=36'h000000000;
			11'h7e5: dataout<=36'h000000000;
			11'h7e6: dataout<=36'h000000000;
			11'h7e7: dataout<=36'h000000000;
			11'h7e8: dataout<=36'h000000000;
			11'h7e9: dataout<=36'h000000000;
			11'h7ea: dataout<=36'h000000000;
			11'h7eb: dataout<=36'h000000000;
			11'h7ec: dataout<=36'h000000000;
			11'h7ed: dataout<=36'h000000000;
			11'h7ee: dataout<=36'h000000000;
			11'h7ef: dataout<=36'h000000000;
			11'h7f0: dataout<=36'h000000000;
			11'h7f1: dataout<=36'h000000000;
			11'h7f2: dataout<=36'h000000000;
			11'h7f3: dataout<=36'h000000000;
			11'h7f4: dataout<=36'h000000000;
			11'h7f5: dataout<=36'h000000000;
			11'h7f6: dataout<=36'h000000000;
			11'h7f7: dataout<=36'h000000000;
			11'h7f8: dataout<=36'h000000000;
			11'h7f9: dataout<=36'h000000000;
			11'h7fa: dataout<=36'h000000000;
			11'h7fb: dataout<=36'h000000000;
			11'h7fc: dataout<=36'h000000000;
			11'h7fd: dataout<=36'h000000000;
			11'h7fe: dataout<=36'h000000000;
			11'h7ff: dataout<=36'h000000000;
		endcase
	end
endmodule

